

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7426, n7427, n7428, n7429, n7430, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625;

  INV_X4 U7527 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X4 U7528 ( .A(n12901), .ZN(n12910) );
  INV_X2 U7529 ( .A(n8620), .ZN(n9342) );
  CLKBUF_X2 U7530 ( .A(n10039), .Z(n9954) );
  INV_X2 U7531 ( .A(n13277), .ZN(n13256) );
  INV_X2 U7532 ( .A(n13345), .ZN(n13105) );
  INV_X1 U7533 ( .A(n9222), .ZN(n9399) );
  NAND2_X1 U7534 ( .A1(n12904), .A2(n12906), .ZN(n12948) );
  INV_X2 U7535 ( .A(n7430), .ZN(n12760) );
  INV_X1 U7536 ( .A(n15252), .ZN(n15223) );
  NAND2_X1 U7537 ( .A1(n8802), .A2(n10468), .ZN(n9321) );
  AND2_X1 U7538 ( .A1(n11366), .A2(n13054), .ZN(n11211) );
  NAND2_X1 U7539 ( .A1(n9966), .A2(n9965), .ZN(n13759) );
  INV_X1 U7540 ( .A(n13779), .ZN(n13421) );
  INV_X1 U7541 ( .A(n13697), .ZN(n7429) );
  INV_X2 U7543 ( .A(n8894), .ZN(n9346) );
  NAND2_X1 U7544 ( .A1(n15351), .A2(n15355), .ZN(n15287) );
  NAND2_X1 U7545 ( .A1(n15969), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10343) );
  OAI21_X1 U7546 ( .B1(n10132), .B2(n8328), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n10218) );
  INV_X2 U7547 ( .A(n10165), .ZN(n10468) );
  OAI21_X1 U7548 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(n16222), .A(n16353), .ZN(
        n16235) );
  NAND2_X1 U7549 ( .A1(n16306), .A2(n7892), .ZN(n16317) );
  NAND4_X2 U7550 ( .A1(n8577), .A2(n8575), .A3(n8576), .A4(n8574), .ZN(n14734)
         );
  INV_X1 U7551 ( .A(n13697), .ZN(n13671) );
  AND2_X1 U7552 ( .A1(n12700), .A2(n12699), .ZN(n7426) );
  NOR2_X1 U7553 ( .A1(n13764), .A2(n12766), .ZN(n12767) );
  AND2_X2 U7554 ( .A1(n9615), .A2(n9616), .ZN(n8365) );
  AND2_X2 U7556 ( .A1(n8345), .A2(n7988), .ZN(n7647) );
  AND2_X2 U7557 ( .A1(n14190), .A2(n10660), .ZN(n14201) );
  NOR2_X2 U7558 ( .A1(n9766), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n9464) );
  NAND2_X2 U7559 ( .A1(n11545), .A2(n11544), .ZN(n12032) );
  NAND2_X2 U7560 ( .A1(n12407), .A2(n12406), .ZN(n15541) );
  NAND2_X2 U7561 ( .A1(n12317), .A2(n8204), .ZN(n12407) );
  INV_X1 U7562 ( .A(n12139), .ZN(n9405) );
  XNOR2_X2 U7563 ( .A(n8529), .B(n8528), .ZN(n12139) );
  NAND2_X2 U7564 ( .A1(n16244), .A2(n16245), .ZN(n16254) );
  OAI22_X2 U7565 ( .A1(n9207), .A2(n8385), .B1(n9208), .B2(n8386), .ZN(n9213)
         );
  INV_X2 U7566 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n10075) );
  OAI21_X2 U7567 ( .B1(n9699), .B2(n9503), .A(n9505), .ZN(n9712) );
  OAI21_X2 U7568 ( .B1(n16298), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n16297), .ZN(
        n16304) );
  XNOR2_X2 U7569 ( .A(n9600), .B(P3_IR_REG_1__SCAN_IN), .ZN(n14155) );
  NAND2_X2 U7570 ( .A1(n9981), .A2(n9980), .ZN(n13741) );
  NAND2_X2 U7571 ( .A1(n9751), .A2(n12839), .ZN(n13964) );
  NAND2_X1 U7572 ( .A1(n13204), .A2(n10468), .ZN(n7428) );
  NAND2_X1 U7573 ( .A1(n13204), .A2(n10468), .ZN(n13290) );
  XNOR2_X2 U7574 ( .A(n8543), .B(n8542), .ZN(n15114) );
  NAND2_X2 U7575 ( .A1(n8541), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8543) );
  XNOR2_X2 U7576 ( .A(n9535), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n9925) );
  OR2_X2 U7577 ( .A1(n7436), .A2(n11536), .ZN(n7443) );
  CLKBUF_X3 U7578 ( .A(n9645), .Z(n7430) );
  NAND2_X1 U7579 ( .A1(n10928), .A2(n10468), .ZN(n9645) );
  INV_X2 U7580 ( .A(n9662), .ZN(n9632) );
  NAND2_X2 U7581 ( .A1(n10219), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10221) );
  NAND2_X2 U7582 ( .A1(n9591), .A2(n9590), .ZN(n10636) );
  NAND2_X2 U7584 ( .A1(n11654), .A2(n11033), .ZN(n9990) );
  AND4_X4 U7585 ( .A1(n9606), .A2(n9605), .A3(n9604), .A4(n7443), .ZN(n11654)
         );
  OAI22_X2 U7586 ( .A1(n10972), .A2(n10973), .B1(n10922), .B2(n10955), .ZN(
        n11223) );
  AOI22_X2 U7587 ( .A1(n11249), .A2(n11248), .B1(n10953), .B2(n10921), .ZN(
        n10972) );
  OAI21_X2 U7588 ( .B1(n9857), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7704) );
  NOR2_X2 U7589 ( .A1(n11224), .A2(n11225), .ZN(n11397) );
  OAI21_X2 U7590 ( .B1(n11223), .B2(n11222), .A(n11221), .ZN(n11224) );
  BUF_X4 U7591 ( .A(n12736), .Z(n7434) );
  NAND2_X2 U7592 ( .A1(n13439), .A2(n14152), .ZN(n12736) );
  AOI21_X2 U7593 ( .B1(n11942), .B2(n9996), .A(n8424), .ZN(n11749) );
  AND2_X2 U7594 ( .A1(n11941), .A2(n9993), .ZN(n9996) );
  NAND2_X2 U7595 ( .A1(n11652), .A2(n9992), .ZN(n11942) );
  INV_X1 U7596 ( .A(n9579), .ZN(n13439) );
  NAND2_X1 U7598 ( .A1(n15694), .A2(n15575), .ZN(n8193) );
  NAND2_X2 U7599 ( .A1(n14081), .A2(n13421), .ZN(n12771) );
  NAND2_X1 U7600 ( .A1(n9962), .A2(n9961), .ZN(n9964) );
  NAND2_X1 U7601 ( .A1(n13903), .A2(n10016), .ZN(n13902) );
  NAND2_X1 U7602 ( .A1(n11811), .A2(n11810), .ZN(n11809) );
  NAND2_X1 U7603 ( .A1(n11940), .A2(n12810), .ZN(n11746) );
  NAND2_X1 U7604 ( .A1(n14168), .A2(n8646), .ZN(n10723) );
  AND4_X1 U7605 ( .A1(n9654), .A2(n9653), .A3(n9652), .A4(n9651), .ZN(n11754)
         );
  INV_X1 U7606 ( .A(n11362), .ZN(n16463) );
  NAND4_X1 U7607 ( .A1(n9668), .A2(n9667), .A3(n9666), .A4(n9665), .ZN(n13605)
         );
  INV_X2 U7608 ( .A(n8016), .ZN(n11689) );
  AND3_X1 U7609 ( .A1(n9661), .A2(n9660), .A3(n9659), .ZN(n11706) );
  NAND4_X1 U7610 ( .A1(n10774), .A2(n10773), .A3(n10772), .A4(n10771), .ZN(
        n15380) );
  CLKBUF_X2 U7611 ( .A(n14884), .Z(n14873) );
  CLKBUF_X2 U7612 ( .A(n14884), .Z(n14986) );
  CLKBUF_X2 U7613 ( .A(n9159), .Z(n9370) );
  OR2_X1 U7614 ( .A1(n8530), .A2(n11319), .ZN(n8598) );
  CLKBUF_X2 U7615 ( .A(n8592), .Z(n9327) );
  INV_X4 U7616 ( .A(n7462), .ZN(n7432) );
  CLKBUF_X2 U7617 ( .A(n10529), .Z(n13282) );
  CLKBUF_X2 U7618 ( .A(n11097), .Z(n7619) );
  INV_X2 U7619 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n14472) );
  MUX2_X1 U7620 ( .A(P3_REG0_REG_28__SCAN_IN), .B(n14071), .S(n16590), .Z(
        n14072) );
  MUX2_X1 U7621 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n14071), .S(n16587), .Z(
        n13991) );
  OR2_X1 U7622 ( .A1(n12919), .A2(n12918), .ZN(n8175) );
  AOI21_X1 U7623 ( .B1(n12917), .B2(n12949), .A(n12916), .ZN(n12919) );
  NOR2_X1 U7624 ( .A1(n15623), .A2(n15624), .ZN(n15622) );
  OAI21_X1 U7625 ( .B1(n13818), .B2(n7983), .A(n7980), .ZN(n13790) );
  INV_X1 U7626 ( .A(n14193), .ZN(n14189) );
  AND2_X1 U7627 ( .A1(n7818), .A2(n7821), .ZN(n15631) );
  NAND2_X1 U7628 ( .A1(n7689), .A2(n7471), .ZN(n15280) );
  NAND2_X1 U7629 ( .A1(n12751), .A2(n12750), .ZN(n13720) );
  NAND2_X1 U7630 ( .A1(n7580), .A2(n7579), .ZN(n13851) );
  AND2_X1 U7631 ( .A1(n14835), .A2(n14834), .ZN(n14837) );
  NAND2_X1 U7632 ( .A1(n8021), .A2(n8019), .ZN(n14652) );
  AND2_X1 U7633 ( .A1(n8995), .A2(n8020), .ZN(n8019) );
  NAND2_X1 U7634 ( .A1(n15041), .A2(n12707), .ZN(n14899) );
  INV_X1 U7635 ( .A(n13759), .ZN(n14076) );
  NAND2_X1 U7636 ( .A1(n7874), .A2(n7873), .ZN(n15724) );
  NAND2_X1 U7637 ( .A1(n7774), .A2(n15741), .ZN(n15735) );
  AOI21_X2 U7638 ( .B1(n13853), .B2(n10026), .A(n8427), .ZN(n13822) );
  NAND2_X1 U7639 ( .A1(n9979), .A2(n9546), .ZN(n12746) );
  NAND2_X1 U7640 ( .A1(n9977), .A2(n9976), .ZN(n9979) );
  NAND2_X1 U7641 ( .A1(n15749), .A2(n15571), .ZN(n15733) );
  INV_X1 U7642 ( .A(n13996), .ZN(n14081) );
  NAND2_X1 U7643 ( .A1(n9963), .A2(n9964), .ZN(n13400) );
  NAND2_X1 U7644 ( .A1(n9964), .A2(n9544), .ZN(n9977) );
  NAND2_X1 U7645 ( .A1(n7702), .A2(n8082), .ZN(n15242) );
  NAND2_X1 U7646 ( .A1(n9938), .A2(n9937), .ZN(n14001) );
  NAND2_X1 U7647 ( .A1(n8237), .A2(n15568), .ZN(n15767) );
  OR2_X1 U7648 ( .A1(n9962), .A2(n9961), .ZN(n9963) );
  OR2_X1 U7649 ( .A1(n12350), .A2(n9644), .ZN(n9938) );
  NAND2_X1 U7650 ( .A1(n9948), .A2(n9947), .ZN(n9949) );
  NOR2_X1 U7651 ( .A1(n13678), .A2(n7642), .ZN(n13679) );
  NAND2_X1 U7652 ( .A1(n8214), .A2(n15655), .ZN(n15632) );
  NAND2_X1 U7653 ( .A1(n15153), .A2(n15154), .ZN(n15353) );
  AND2_X1 U7654 ( .A1(n15148), .A2(n15147), .ZN(n15153) );
  AND2_X1 U7655 ( .A1(n12869), .A2(n12870), .ZN(n13876) );
  NAND2_X1 U7656 ( .A1(n12362), .A2(n12361), .ZN(n12516) );
  OR2_X1 U7657 ( .A1(n12436), .A2(n12437), .ZN(n7909) );
  XNOR2_X1 U7658 ( .A(n12485), .B(n12486), .ZN(n12436) );
  OR2_X1 U7659 ( .A1(n9046), .A2(n9045), .ZN(n9048) );
  NAND2_X1 U7660 ( .A1(n11964), .A2(n11963), .ZN(n12020) );
  AND2_X1 U7661 ( .A1(n12435), .A2(n12441), .ZN(n12485) );
  NAND2_X1 U7662 ( .A1(n16293), .A2(n16292), .ZN(n16295) );
  NAND2_X1 U7663 ( .A1(n12634), .A2(n8886), .ZN(n8897) );
  NAND2_X1 U7664 ( .A1(n9945), .A2(n9944), .ZN(n13795) );
  AND2_X1 U7665 ( .A1(n9862), .A2(n9861), .ZN(n13884) );
  AND2_X1 U7666 ( .A1(n12375), .A2(n12374), .ZN(n12377) );
  OAI21_X1 U7667 ( .B1(n11809), .B2(n7564), .A(n8234), .ZN(n11966) );
  NAND2_X1 U7668 ( .A1(n11415), .A2(n11414), .ZN(n11612) );
  OR2_X1 U7669 ( .A1(n12501), .A2(n7554), .ZN(n7640) );
  NAND2_X1 U7670 ( .A1(n11375), .A2(n8748), .ZN(n11460) );
  NAND2_X1 U7671 ( .A1(n12243), .A2(n10003), .ZN(n12291) );
  NAND2_X1 U7672 ( .A1(n9806), .A2(n9517), .ZN(n9819) );
  AND2_X1 U7673 ( .A1(n12839), .A2(n12840), .ZN(n12936) );
  OAI21_X1 U7674 ( .B1(n11360), .B2(n13048), .A(n13050), .ZN(n11055) );
  OAI211_X1 U7675 ( .C1(n11349), .C2(n8070), .A(n11351), .B(n7772), .ZN(n11549) );
  NAND2_X1 U7676 ( .A1(n7884), .A2(n7883), .ZN(n16245) );
  NAND2_X1 U7677 ( .A1(n11649), .A2(n9619), .ZN(n12792) );
  INV_X2 U7678 ( .A(n16622), .ZN(n7433) );
  AND3_X1 U7679 ( .A1(n9735), .A2(n9734), .A3(n9733), .ZN(n12546) );
  OAI21_X1 U7680 ( .B1(n11740), .B2(n11739), .A(n11738), .ZN(n11769) );
  INV_X1 U7681 ( .A(n16239), .ZN(n7884) );
  NAND2_X1 U7682 ( .A1(n9730), .A2(n9729), .ZN(n9728) );
  NAND2_X1 U7683 ( .A1(n8206), .A2(n16452), .ZN(n11363) );
  NAND2_X1 U7684 ( .A1(n8734), .A2(n8733), .ZN(n12095) );
  NAND2_X1 U7685 ( .A1(n9714), .A2(n9507), .ZN(n9730) );
  AND2_X2 U7686 ( .A1(n15589), .A2(n16395), .ZN(n16605) );
  NAND2_X1 U7687 ( .A1(n11292), .A2(n11291), .ZN(n16526) );
  NAND2_X1 U7688 ( .A1(n11030), .A2(n11029), .ZN(n11499) );
  AND3_X1 U7689 ( .A1(n9691), .A2(n9690), .A3(n9689), .ZN(n13445) );
  AND3_X1 U7690 ( .A1(n9674), .A2(n9673), .A3(n9672), .ZN(n12814) );
  NAND4_X1 U7691 ( .A1(n9727), .A2(n9726), .A3(n9725), .A4(n9724), .ZN(n12832)
         );
  NAND2_X1 U7692 ( .A1(n8711), .A2(n8710), .ZN(n8713) );
  AND4_X1 U7693 ( .A1(n9636), .A2(n9635), .A3(n9634), .A4(n9633), .ZN(n9646)
         );
  NAND4_X1 U7694 ( .A1(n9611), .A2(n9610), .A3(n9609), .A4(n9608), .ZN(n11194)
         );
  NAND2_X1 U7695 ( .A1(n7577), .A2(n7576), .ZN(n9684) );
  NOR2_X1 U7696 ( .A1(n16205), .A2(n16206), .ZN(n16220) );
  INV_X1 U7697 ( .A(n9168), .ZN(n9222) );
  INV_X2 U7698 ( .A(n8598), .ZN(n14190) );
  INV_X2 U7699 ( .A(n9662), .ZN(n7437) );
  OAI211_X1 U7700 ( .C1(SI_2_), .C2(n9645), .A(n9618), .B(n9617), .ZN(n12798)
         );
  AND4_X1 U7701 ( .A1(n10536), .A2(n10535), .A3(n10534), .A4(n10533), .ZN(
        n10878) );
  AOI21_X1 U7702 ( .B1(n11228), .B2(n11227), .A(n7615), .ZN(n11383) );
  NAND4_X1 U7703 ( .A1(n8596), .A2(n8593), .A3(n8594), .A4(n8595), .ZN(n14737)
         );
  NAND4_X2 U7704 ( .A1(n8580), .A2(n7473), .A3(n8581), .A4(n8582), .ZN(n14735)
         );
  OR2_X1 U7705 ( .A1(n9752), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9781) );
  INV_X1 U7706 ( .A(n12739), .ZN(n7435) );
  INV_X2 U7707 ( .A(n9644), .ZN(n12759) );
  AND2_X2 U7708 ( .A1(n12988), .A2(n12987), .ZN(n13345) );
  OAI22_X1 U7709 ( .A1(n10974), .A2(n10944), .B1(n10943), .B2(n10978), .ZN(
        n11228) );
  NAND2_X1 U7710 ( .A1(n9579), .A2(n14152), .ZN(n12739) );
  INV_X1 U7711 ( .A(n10928), .ZN(n9768) );
  NAND2_X2 U7712 ( .A1(n8545), .A2(n12730), .ZN(n8620) );
  AND2_X2 U7713 ( .A1(n12730), .A2(n15114), .ZN(n8894) );
  AND2_X1 U7714 ( .A1(n9155), .A2(n9405), .ZN(n11319) );
  INV_X2 U7715 ( .A(n12973), .ZN(n13289) );
  NAND2_X1 U7716 ( .A1(n13027), .A2(n10410), .ZN(n7462) );
  NAND2_X2 U7717 ( .A1(n9578), .A2(n14144), .ZN(n14152) );
  NOR2_X1 U7718 ( .A1(n9824), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n9826) );
  NAND2_X1 U7719 ( .A1(n9554), .A2(n9575), .ZN(n12732) );
  INV_X1 U7720 ( .A(n10036), .ZN(n13697) );
  CLKBUF_X1 U7721 ( .A(n9154), .Z(n11851) );
  MUX2_X1 U7722 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9553), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n9554) );
  XNOR2_X1 U7723 ( .A(n10337), .B(n8109), .ZN(n12993) );
  AND2_X1 U7724 ( .A1(n9643), .A2(n9642), .ZN(n10953) );
  XNOR2_X1 U7725 ( .A(n10347), .B(n10346), .ZN(n15979) );
  NAND2_X1 U7726 ( .A1(n8508), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8510) );
  OAI21_X1 U7727 ( .B1(n8889), .B2(n8521), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8524) );
  NAND2_X1 U7728 ( .A1(n8080), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8079) );
  XNOR2_X1 U7729 ( .A(n10218), .B(n10217), .ZN(n13373) );
  OAI21_X1 U7730 ( .B1(n8461), .B2(SI_9_), .A(n8463), .ZN(n8730) );
  OR2_X1 U7731 ( .A1(n10345), .A2(n10344), .ZN(n10347) );
  AND2_X1 U7732 ( .A1(n9547), .A2(n7989), .ZN(n8346) );
  NAND2_X1 U7733 ( .A1(n10131), .A2(n10220), .ZN(n8328) );
  NOR2_X1 U7734 ( .A1(n8367), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8364) );
  AND2_X1 U7735 ( .A1(n10170), .A2(n14579), .ZN(n10166) );
  AND4_X1 U7736 ( .A1(n9457), .A2(n9456), .A3(n9685), .A4(n9731), .ZN(n9458)
         );
  AND3_X1 U7737 ( .A1(n10130), .A2(n10137), .A3(n10129), .ZN(n10131) );
  NOR2_X1 U7738 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n16167), .ZN(n16172) );
  AND4_X1 U7739 ( .A1(n10111), .A2(n10110), .A3(n10109), .A4(n14380), .ZN(
        n7685) );
  AND3_X1 U7740 ( .A1(n10114), .A2(n10113), .A3(n10112), .ZN(n10249) );
  INV_X4 U7741 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U7742 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n10110) );
  NOR2_X1 U7743 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n10109) );
  INV_X1 U7744 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n14380) );
  INV_X1 U7745 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10493) );
  NOR2_X1 U7746 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n10113) );
  NOR2_X1 U7747 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n10112) );
  INV_X1 U7748 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8906) );
  NOR2_X1 U7749 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8497) );
  INV_X1 U7750 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8515) );
  INV_X1 U7751 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9731) );
  INV_X1 U7752 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9685) );
  INV_X1 U7753 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9548) );
  NOR2_X1 U7754 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n9456) );
  NOR2_X1 U7755 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n9457) );
  INV_X1 U7756 ( .A(n14170), .ZN(n11990) );
  AOI21_X2 U7757 ( .B1(n11681), .B2(n11680), .A(n11679), .ZN(n11740) );
  BUF_X4 U7758 ( .A(n12739), .Z(n7436) );
  OAI21_X4 U7759 ( .B1(n9917), .B2(n9916), .A(n9534), .ZN(n9535) );
  OR2_X1 U7760 ( .A1(n7434), .A2(n9599), .ZN(n9604) );
  OAI21_X2 U7761 ( .B1(n15541), .B2(n7869), .A(n7866), .ZN(n15763) );
  OAI222_X1 U7762 ( .A1(P1_U3086), .A2(n15976), .B1(n15990), .B2(n15975), .C1(
        n15974), .C2(n15987), .ZN(P1_U3325) );
  INV_X2 U7763 ( .A(n13025), .ZN(n7601) );
  OAI21_X2 U7764 ( .B1(n9762), .B2(n8166), .A(n8162), .ZN(n9789) );
  NAND2_X2 U7765 ( .A1(n9758), .A2(n9759), .ZN(n9762) );
  INV_X1 U7766 ( .A(n8178), .ZN(n8211) );
  OAI222_X1 U7767 ( .A1(n13439), .A2(P3_U3151), .B1(n14150), .B2(n13438), .C1(
        n14154), .C2(n13437), .ZN(P3_U3265) );
  MUX2_X2 U7768 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9576), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n9578) );
  MUX2_X2 U7769 ( .A(n10105), .B(n10104), .S(n16590), .Z(n10108) );
  MUX2_X2 U7770 ( .A(n10087), .B(n10104), .S(n16587), .Z(n10091) );
  AOI21_X2 U7771 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(n16256), .A(n16255), .ZN(
        n16268) );
  OAI222_X1 U7772 ( .A1(n14154), .A2(n14153), .B1(P3_U3151), .B2(n14152), .C1(
        n14151), .C2(n14150), .ZN(P3_U3266) );
  INV_X1 U7773 ( .A(n14152), .ZN(n9580) );
  XNOR2_X1 U7774 ( .A(n12734), .B(n12903), .ZN(n13723) );
  NAND2_X2 U7775 ( .A1(n13838), .A2(n13401), .ZN(n13818) );
  AND2_X4 U7776 ( .A1(n7860), .A2(n7858), .ZN(n16434) );
  INV_X1 U7777 ( .A(n8956), .ZN(n8957) );
  NAND2_X1 U7778 ( .A1(n8935), .A2(n8938), .ZN(n8285) );
  AOI21_X1 U7779 ( .B1(n8274), .B2(n8275), .A(n8272), .ZN(n8271) );
  INV_X1 U7780 ( .A(n8849), .ZN(n8272) );
  NAND2_X1 U7781 ( .A1(n7478), .A2(n10027), .ZN(n8000) );
  INV_X1 U7782 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9552) );
  OR2_X1 U7783 ( .A1(n11346), .A2(n11345), .ZN(n11349) );
  OAI21_X1 U7784 ( .B1(n9355), .B2(n9354), .A(n9301), .ZN(n9338) );
  NAND2_X1 U7785 ( .A1(n8474), .A2(n8473), .ZN(n8812) );
  NAND2_X1 U7786 ( .A1(n7810), .A2(n7809), .ZN(n15596) );
  XNOR2_X1 U7787 ( .A(n15840), .B(n15370), .ZN(n15624) );
  NAND2_X1 U7788 ( .A1(n7878), .A2(n7875), .ZN(n15647) );
  NOR2_X1 U7789 ( .A1(n15650), .A2(n8183), .ZN(n7875) );
  NAND2_X1 U7790 ( .A1(n11806), .A2(n11584), .ZN(n11589) );
  NAND2_X1 U7791 ( .A1(n13204), .A2(n10165), .ZN(n12973) );
  NAND2_X2 U7792 ( .A1(n13373), .A2(n15982), .ZN(n13204) );
  NAND2_X1 U7793 ( .A1(n9163), .A2(n9162), .ZN(n7827) );
  OR2_X1 U7794 ( .A1(n9194), .A2(n7853), .ZN(n7852) );
  INV_X1 U7795 ( .A(n9193), .ZN(n7853) );
  NAND2_X1 U7796 ( .A1(n9219), .A2(n8393), .ZN(n8392) );
  INV_X1 U7797 ( .A(n9220), .ZN(n8393) );
  NAND2_X1 U7798 ( .A1(n7574), .A2(n7573), .ZN(n7572) );
  NOR2_X1 U7799 ( .A1(n12777), .A2(n12901), .ZN(n7573) );
  NAND2_X1 U7800 ( .A1(n12897), .A2(n12778), .ZN(n7574) );
  NAND2_X1 U7801 ( .A1(n7591), .A2(n9415), .ZN(n9383) );
  NAND2_X1 U7802 ( .A1(n7672), .A2(n7494), .ZN(n13298) );
  INV_X1 U7803 ( .A(n8490), .ZN(n7924) );
  AOI21_X1 U7804 ( .B1(n8271), .B2(n8273), .A(n7512), .ZN(n7942) );
  INV_X1 U7805 ( .A(n8274), .ZN(n8273) );
  INV_X1 U7806 ( .A(n13953), .ZN(n13376) );
  AND2_X1 U7807 ( .A1(n7525), .A2(n7446), .ZN(n8376) );
  OR2_X1 U7808 ( .A1(n14020), .A2(n13855), .ZN(n13402) );
  NAND2_X1 U7809 ( .A1(n13766), .A2(n10031), .ZN(n8009) );
  OR2_X1 U7810 ( .A1(n13811), .A2(n13824), .ZN(n12893) );
  AOI21_X1 U7811 ( .B1(n7999), .B2(n7997), .A(n7499), .ZN(n7996) );
  INV_X1 U7812 ( .A(n10027), .ZN(n7997) );
  NOR2_X1 U7813 ( .A1(n10020), .A2(n7476), .ZN(n8015) );
  INV_X1 U7814 ( .A(n12963), .ZN(n9480) );
  OR2_X1 U7815 ( .A1(n9555), .A2(n14143), .ZN(n9557) );
  AND3_X1 U7816 ( .A1(n9467), .A2(n9466), .A3(n9465), .ZN(n9547) );
  NAND2_X1 U7817 ( .A1(n10205), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9502) );
  OR2_X1 U7818 ( .A1(n9290), .A2(n9289), .ZN(n7612) );
  AND2_X1 U7819 ( .A1(n9396), .A2(n9375), .ZN(n9376) );
  INV_X1 U7820 ( .A(n9293), .ZN(n7847) );
  XNOR2_X1 U7821 ( .A(n14804), .B(n14807), .ZN(n9415) );
  INV_X1 U7822 ( .A(n12730), .ZN(n8544) );
  INV_X1 U7823 ( .A(n15114), .ZN(n8545) );
  OR2_X1 U7824 ( .A1(n15011), .A2(n9416), .ZN(n12690) );
  NOR2_X1 U7825 ( .A1(n8057), .A2(n7503), .ZN(n8056) );
  INV_X1 U7826 ( .A(n12685), .ZN(n8057) );
  NAND2_X1 U7827 ( .A1(n9030), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9054) );
  OR2_X1 U7828 ( .A1(n12642), .A2(n7762), .ZN(n7761) );
  NOR2_X1 U7829 ( .A1(n12590), .A2(n8055), .ZN(n8054) );
  INV_X1 U7830 ( .A(n12567), .ZN(n8055) );
  AND2_X1 U7831 ( .A1(n10870), .A2(n13028), .ZN(n15221) );
  INV_X1 U7832 ( .A(n15976), .ZN(n10348) );
  NOR2_X1 U7833 ( .A1(n8231), .A2(n7873), .ZN(n8230) );
  INV_X1 U7834 ( .A(n15576), .ZN(n8231) );
  INV_X1 U7835 ( .A(n8181), .ZN(n8180) );
  OAI21_X1 U7836 ( .B1(n15816), .B2(n8182), .A(n15544), .ZN(n8181) );
  INV_X1 U7837 ( .A(n8218), .ZN(n8217) );
  OAI21_X1 U7838 ( .B1(n12003), .B2(n8219), .A(n12408), .ZN(n8218) );
  NAND2_X1 U7839 ( .A1(n8259), .A2(n8258), .ZN(n9355) );
  AOI21_X1 U7840 ( .B1(n8261), .B2(n8263), .A(n7569), .ZN(n8258) );
  NAND2_X1 U7841 ( .A1(n9024), .A2(n9023), .ZN(n9046) );
  NAND2_X1 U7842 ( .A1(n7925), .A2(n8490), .ZN(n8936) );
  NAND2_X1 U7843 ( .A1(n7926), .A2(n8257), .ZN(n7925) );
  AND2_X1 U7844 ( .A1(n8487), .A2(n7927), .ZN(n7926) );
  XNOR2_X1 U7845 ( .A(n8488), .B(SI_19_), .ZN(n8551) );
  NAND2_X1 U7846 ( .A1(n7797), .A2(n7794), .ZN(n8485) );
  OR2_X1 U7847 ( .A1(n7800), .A2(n7799), .ZN(n7797) );
  OAI21_X1 U7848 ( .B1(n8868), .B2(n7798), .A(n14425), .ZN(n7795) );
  XNOR2_X1 U7849 ( .A(n8483), .B(SI_17_), .ZN(n8887) );
  OR2_X1 U7850 ( .A1(n8868), .A2(n8867), .ZN(n8870) );
  NAND2_X1 U7851 ( .A1(n7786), .A2(n7787), .ZN(n8789) );
  AND2_X1 U7852 ( .A1(n7788), .A2(n7928), .ZN(n7787) );
  AOI21_X1 U7853 ( .B1(n8749), .B2(n7930), .A(n7516), .ZN(n7928) );
  NAND2_X1 U7854 ( .A1(n8650), .A2(n7741), .ZN(n7740) );
  INV_X1 U7855 ( .A(n8445), .ZN(n7741) );
  AND2_X1 U7856 ( .A1(n8650), .A2(n8443), .ZN(n7610) );
  INV_X1 U7857 ( .A(n8568), .ZN(n7944) );
  INV_X1 U7858 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n16217) );
  NAND2_X1 U7859 ( .A1(n12457), .A2(n12456), .ZN(n7720) );
  NAND2_X1 U7860 ( .A1(n12157), .A2(n8333), .ZN(n12387) );
  NOR2_X1 U7861 ( .A1(n12160), .A2(n8334), .ZN(n8333) );
  INV_X1 U7862 ( .A(n12156), .ZN(n8334) );
  NOR2_X1 U7863 ( .A1(n11728), .A2(n11727), .ZN(n11766) );
  NAND2_X1 U7864 ( .A1(n7899), .A2(n11897), .ZN(n12435) );
  NAND2_X1 U7865 ( .A1(n7737), .A2(n7736), .ZN(n13609) );
  INV_X1 U7866 ( .A(n12490), .ZN(n7736) );
  XNOR2_X1 U7867 ( .A(n13811), .B(n13824), .ZN(n13808) );
  NAND2_X1 U7868 ( .A1(n13889), .A2(n10018), .ZN(n13875) );
  OAI21_X1 U7869 ( .B1(n12291), .B2(n12462), .A(n12544), .ZN(n10005) );
  NAND2_X1 U7870 ( .A1(n9480), .A2(n11442), .ZN(n16580) );
  XNOR2_X1 U7871 ( .A(n10058), .B(P3_IR_REG_26__SCAN_IN), .ZN(n10079) );
  OR2_X1 U7872 ( .A1(n9473), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n10074) );
  NAND2_X1 U7873 ( .A1(n9826), .A2(n9462), .ZN(n9857) );
  NAND2_X1 U7874 ( .A1(n8167), .A2(n8168), .ZN(n9773) );
  CLKBUF_X1 U7875 ( .A(n9765), .Z(n9766) );
  CLKBUF_X1 U7876 ( .A(n9156), .Z(n8519) );
  NAND2_X1 U7877 ( .A1(n8074), .A2(n12690), .ZN(n7773) );
  NOR2_X1 U7878 ( .A1(n14844), .A2(n15011), .ZN(n14824) );
  AND2_X1 U7879 ( .A1(n9140), .A2(n9079), .ZN(n14846) );
  NAND2_X1 U7880 ( .A1(n14939), .A2(n14938), .ZN(n7771) );
  OAI21_X1 U7881 ( .B1(n14964), .B2(n12677), .A(n12676), .ZN(n14946) );
  NAND2_X1 U7882 ( .A1(n14968), .A2(n12701), .ZN(n14945) );
  AND2_X1 U7883 ( .A1(n12268), .A2(n9419), .ZN(n12194) );
  NAND2_X1 U7884 ( .A1(n11549), .A2(n12024), .ZN(n11550) );
  INV_X1 U7885 ( .A(n14884), .ZN(n14930) );
  XNOR2_X1 U7886 ( .A(n14170), .B(n14733), .ZN(n10815) );
  XNOR2_X1 U7887 ( .A(n8524), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9154) );
  INV_X1 U7888 ( .A(n8097), .ZN(n8096) );
  OAI21_X1 U7889 ( .B1(n15343), .B2(n8101), .A(n15341), .ZN(n8097) );
  OR2_X1 U7890 ( .A1(n10876), .A2(n15223), .ZN(n10521) );
  NAND2_X1 U7891 ( .A1(n8114), .A2(n7485), .ZN(n15269) );
  OR2_X1 U7892 ( .A1(n15211), .A2(n15210), .ZN(n7695) );
  OR2_X1 U7893 ( .A1(n15303), .A2(n7696), .ZN(n7694) );
  OAI21_X1 U7894 ( .B1(n13363), .B2(n7663), .A(n13364), .ZN(n7662) );
  NAND2_X1 U7895 ( .A1(n7665), .A2(n7664), .ZN(n7663) );
  NOR2_X1 U7896 ( .A1(n13361), .A2(n13360), .ZN(n7664) );
  NAND2_X1 U7897 ( .A1(n10348), .A2(n10350), .ZN(n10529) );
  NOR2_X1 U7898 ( .A1(n13305), .A2(n8209), .ZN(n8207) );
  NOR2_X1 U7899 ( .A1(n15622), .A2(n7549), .ZN(n15602) );
  NAND2_X1 U7900 ( .A1(n15628), .A2(n8428), .ZN(n15623) );
  OR2_X1 U7901 ( .A1(n15580), .A2(n15653), .ZN(n8428) );
  NAND2_X1 U7902 ( .A1(n15635), .A2(n15621), .ZN(n15615) );
  INV_X1 U7903 ( .A(n15867), .ZN(n15686) );
  NAND2_X1 U7904 ( .A1(n15888), .A2(n15551), .ZN(n15725) );
  NOR2_X1 U7905 ( .A1(n15764), .A2(n8238), .ZN(n8237) );
  INV_X1 U7906 ( .A(n15567), .ZN(n8238) );
  NOR2_X1 U7907 ( .A1(n13329), .A2(n8205), .ZN(n8204) );
  INV_X1 U7908 ( .A(n12316), .ZN(n8205) );
  NAND2_X1 U7909 ( .A1(n12021), .A2(n13328), .ZN(n12317) );
  NOR2_X1 U7910 ( .A1(n13324), .A2(n8187), .ZN(n8186) );
  INV_X1 U7911 ( .A(n11860), .ZN(n8187) );
  NAND2_X1 U7912 ( .A1(n11589), .A2(n11588), .ZN(n11861) );
  NAND2_X1 U7913 ( .A1(n8222), .A2(n8220), .ZN(n11811) );
  OR2_X1 U7914 ( .A1(n8224), .A2(n8221), .ZN(n8220) );
  INV_X1 U7915 ( .A(n11591), .ZN(n8221) );
  NOR2_X1 U7916 ( .A1(n13320), .A2(n8185), .ZN(n8184) );
  INV_X1 U7917 ( .A(n11561), .ZN(n8185) );
  NAND2_X1 U7918 ( .A1(n10877), .A2(n13042), .ZN(n11360) );
  AND2_X1 U7919 ( .A1(n12983), .A2(n12999), .ZN(n16386) );
  AOI21_X1 U7920 ( .B1(n15104), .B2(n13289), .A(n12967), .ZN(n15823) );
  INV_X1 U7921 ( .A(n15621), .ZN(n15840) );
  NOR2_X1 U7922 ( .A1(n15687), .A2(n8192), .ZN(n8191) );
  INV_X1 U7923 ( .A(n15555), .ZN(n8192) );
  AND2_X1 U7924 ( .A1(n10410), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10179) );
  NAND2_X1 U7925 ( .A1(n8326), .A2(n10131), .ZN(n10219) );
  INV_X1 U7926 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n14606) );
  NAND2_X1 U7927 ( .A1(n8270), .A2(n8274), .ZN(n8850) );
  NAND2_X1 U7928 ( .A1(n8812), .A2(n8276), .ZN(n8270) );
  AND2_X1 U7929 ( .A1(n14196), .A2(n14197), .ZN(n7632) );
  NAND2_X1 U7930 ( .A1(n8073), .A2(n7609), .ZN(n7608) );
  INV_X1 U7931 ( .A(n14823), .ZN(n7609) );
  XNOR2_X1 U7932 ( .A(n15583), .B(n15582), .ZN(n15832) );
  AND2_X1 U7933 ( .A1(n8242), .A2(n8241), .ZN(n15842) );
  AOI21_X1 U7934 ( .B1(n15613), .B2(n15789), .A(n7546), .ZN(n8241) );
  NAND2_X1 U7935 ( .A1(n8243), .A2(n16458), .ZN(n8242) );
  OAI21_X1 U7936 ( .B1(n7827), .B2(n7826), .A(n7825), .ZN(n7824) );
  AND2_X1 U7937 ( .A1(n9165), .A2(n9164), .ZN(n7826) );
  NAND2_X1 U7938 ( .A1(n9222), .A2(n14734), .ZN(n9169) );
  NAND2_X1 U7939 ( .A1(n8291), .A2(n7472), .ZN(n7656) );
  NAND2_X1 U7940 ( .A1(n13084), .A2(n7659), .ZN(n7658) );
  AND2_X1 U7941 ( .A1(n7535), .A2(n7657), .ZN(n7655) );
  NAND2_X1 U7942 ( .A1(n13083), .A2(n13085), .ZN(n7657) );
  INV_X1 U7943 ( .A(n7541), .ZN(n7833) );
  NAND2_X1 U7944 ( .A1(n8387), .A2(n7541), .ZN(n7831) );
  NAND2_X1 U7945 ( .A1(n13099), .A2(n13101), .ZN(n8297) );
  AOI21_X1 U7946 ( .B1(n9200), .B2(n9199), .A(n9198), .ZN(n9202) );
  INV_X1 U7947 ( .A(n9227), .ZN(n7623) );
  OR2_X1 U7948 ( .A1(n9215), .A2(n9214), .ZN(n9221) );
  NAND2_X1 U7949 ( .A1(n8390), .A2(n9227), .ZN(n8389) );
  INV_X1 U7950 ( .A(n8392), .ZN(n8390) );
  NAND2_X1 U7951 ( .A1(n8395), .A2(n9227), .ZN(n8391) );
  AOI21_X1 U7952 ( .B1(n9235), .B2(n8407), .A(n8405), .ZN(n8404) );
  NAND2_X1 U7953 ( .A1(n8406), .A2(n9241), .ZN(n8405) );
  NAND2_X1 U7954 ( .A1(n8410), .A2(n8407), .ZN(n8406) );
  OR2_X1 U7955 ( .A1(n8320), .A2(n13165), .ZN(n8318) );
  NAND2_X1 U7956 ( .A1(n7680), .A2(n7508), .ZN(n7679) );
  NAND2_X1 U7957 ( .A1(n7681), .A2(n8319), .ZN(n7680) );
  INV_X1 U7958 ( .A(n8319), .ZN(n7683) );
  NAND2_X1 U7959 ( .A1(n13194), .A2(n8309), .ZN(n8306) );
  NOR2_X1 U7960 ( .A1(n7452), .A2(n7839), .ZN(n7837) );
  NAND2_X1 U7961 ( .A1(n7677), .A2(n13241), .ZN(n7675) );
  NAND2_X1 U7962 ( .A1(n13254), .A2(n8313), .ZN(n8310) );
  NAND2_X1 U7963 ( .A1(n13294), .A2(n13293), .ZN(n8324) );
  INV_X1 U7964 ( .A(n13274), .ZN(n8325) );
  AND2_X1 U7965 ( .A1(n8358), .A2(n8356), .ZN(n8355) );
  OR2_X1 U7966 ( .A1(n13694), .A2(n12789), .ZN(n11025) );
  NAND2_X1 U7967 ( .A1(n7578), .A2(n9994), .ZN(n11943) );
  AND2_X1 U7968 ( .A1(n9052), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n9076) );
  NAND2_X1 U7969 ( .A1(n15580), .A2(n15614), .ZN(n7822) );
  AND2_X1 U7970 ( .A1(n12984), .A2(n12993), .ZN(n13027) );
  NAND2_X1 U7971 ( .A1(n15519), .A2(n12993), .ZN(n12980) );
  NOR2_X1 U7972 ( .A1(n8996), .A2(n8256), .ZN(n8255) );
  AOI21_X1 U7973 ( .B1(n8462), .B2(n7793), .A(n7792), .ZN(n7791) );
  INV_X1 U7974 ( .A(n8463), .ZN(n7792) );
  INV_X1 U7975 ( .A(n8460), .ZN(n7793) );
  NAND2_X1 U7976 ( .A1(n8461), .A2(SI_9_), .ZN(n8463) );
  INV_X1 U7977 ( .A(SI_3_), .ZN(n7753) );
  NOR2_X1 U7978 ( .A1(n8608), .A2(n7758), .ZN(n8612) );
  AND2_X1 U7979 ( .A1(n8568), .A2(n10150), .ZN(n7758) );
  OR2_X1 U7980 ( .A1(n12548), .A2(n8344), .ZN(n8343) );
  INV_X1 U7981 ( .A(n12615), .ZN(n8344) );
  AND2_X1 U7982 ( .A1(n7448), .A2(n7715), .ZN(n7714) );
  NAND2_X1 U7983 ( .A1(n7718), .A2(n7716), .ZN(n7715) );
  INV_X1 U7984 ( .A(n12456), .ZN(n7716) );
  NAND2_X1 U7985 ( .A1(n7714), .A2(n7717), .ZN(n7713) );
  INV_X1 U7986 ( .A(n7718), .ZN(n7717) );
  INV_X1 U7987 ( .A(n13586), .ZN(n8361) );
  AOI21_X1 U7988 ( .B1(n8355), .B2(n8353), .A(n13594), .ZN(n8350) );
  AOI21_X1 U7989 ( .B1(n8353), .B2(n8358), .A(n8356), .ZN(n8352) );
  INV_X1 U7990 ( .A(n8355), .ZN(n8351) );
  NOR2_X1 U7991 ( .A1(n8426), .A2(n7719), .ZN(n7718) );
  INV_X1 U7992 ( .A(n12459), .ZN(n7719) );
  NAND2_X1 U7993 ( .A1(n8374), .A2(n8372), .ZN(n8371) );
  INV_X1 U7994 ( .A(n13388), .ZN(n8372) );
  OR2_X1 U7995 ( .A1(n13389), .A2(n8373), .ZN(n8369) );
  INV_X1 U7996 ( .A(n8374), .ZN(n8373) );
  NAND2_X1 U7997 ( .A1(n7575), .A2(n7572), .ZN(n12900) );
  NAND2_X1 U7998 ( .A1(n12903), .A2(n12902), .ZN(n7628) );
  AND2_X1 U7999 ( .A1(n10012), .A2(n10011), .ZN(n8010) );
  NAND2_X1 U8000 ( .A1(n8009), .A2(n7496), .ZN(n13748) );
  OR2_X1 U8001 ( .A1(n13801), .A2(n13807), .ZN(n12781) );
  NOR2_X1 U8002 ( .A1(n13808), .A2(n7985), .ZN(n7984) );
  INV_X1 U8003 ( .A(n9915), .ZN(n7985) );
  INV_X1 U8004 ( .A(n7972), .ZN(n7971) );
  OAI21_X1 U8005 ( .B1(n13876), .B2(n7973), .A(n13864), .ZN(n7972) );
  OR2_X1 U8006 ( .A1(n14023), .A2(n13867), .ZN(n12879) );
  NOR2_X1 U8007 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_28__SCAN_IN), .ZN(
        n8381) );
  NAND2_X1 U8008 ( .A1(n9536), .A2(n9539), .ZN(n8147) );
  INV_X1 U8009 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n9550) );
  INV_X1 U8010 ( .A(n9853), .ZN(n8160) );
  NOR2_X1 U8011 ( .A1(n9838), .A2(n8159), .ZN(n8158) );
  INV_X1 U8012 ( .A(n9520), .ZN(n8159) );
  INV_X1 U8013 ( .A(n9291), .ZN(n7611) );
  NAND2_X1 U8014 ( .A1(n8398), .A2(n8399), .ZN(n9288) );
  AOI21_X1 U8015 ( .B1(n8398), .B2(n8396), .A(n9287), .ZN(n7855) );
  INV_X1 U8016 ( .A(n9374), .ZN(n7850) );
  INV_X1 U8017 ( .A(n9373), .ZN(n7849) );
  NOR2_X1 U8018 ( .A1(n9388), .A2(n9369), .ZN(n9396) );
  NAND2_X1 U8019 ( .A1(n12714), .A2(n12713), .ZN(n8136) );
  INV_X1 U8020 ( .A(n8056), .ZN(n7749) );
  OR2_X1 U8021 ( .A1(n7953), .A2(n14860), .ZN(n12711) );
  INV_X1 U8022 ( .A(n12708), .ZN(n8127) );
  INV_X1 U8023 ( .A(n12673), .ZN(n7762) );
  INV_X1 U8024 ( .A(n12194), .ZN(n7769) );
  AOI21_X1 U8025 ( .B1(n12194), .B2(n7768), .A(n7767), .ZN(n7766) );
  INV_X1 U8026 ( .A(n12268), .ZN(n7767) );
  INV_X1 U8027 ( .A(n12191), .ZN(n7768) );
  AND2_X1 U8028 ( .A1(n12073), .A2(n12071), .ZN(n8146) );
  OR2_X1 U8029 ( .A1(n12151), .A2(n8069), .ZN(n8067) );
  OR2_X1 U8030 ( .A1(n12142), .A2(n8068), .ZN(n8066) );
  AND2_X1 U8031 ( .A1(n12151), .A2(n8069), .ZN(n8068) );
  NAND2_X1 U8032 ( .A1(n8533), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8777) );
  INV_X1 U8033 ( .A(n8756), .ZN(n8533) );
  NAND2_X1 U8034 ( .A1(n12033), .A2(n11546), .ZN(n8141) );
  INV_X1 U8035 ( .A(n11546), .ZN(n8138) );
  INV_X1 U8036 ( .A(n11342), .ZN(n8123) );
  INV_X1 U8037 ( .A(n7466), .ZN(n8121) );
  NOR2_X1 U8038 ( .A1(n7456), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n8049) );
  OR2_X1 U8039 ( .A1(n8732), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8790) );
  INV_X1 U8040 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8493) );
  NOR2_X1 U8041 ( .A1(n7471), .A2(n7691), .ZN(n7690) );
  OAI21_X1 U8042 ( .B1(n13298), .B2(n13297), .A(n13296), .ZN(n13299) );
  INV_X1 U8043 ( .A(n15837), .ZN(n8210) );
  AND2_X1 U8044 ( .A1(n8180), .A2(n7871), .ZN(n7870) );
  NAND2_X1 U8045 ( .A1(n15559), .A2(n7872), .ZN(n7871) );
  INV_X1 U8046 ( .A(n15543), .ZN(n8182) );
  NAND2_X1 U8047 ( .A1(n7870), .A2(n7868), .ZN(n7867) );
  INV_X1 U8048 ( .A(n7872), .ZN(n7868) );
  OR2_X1 U8049 ( .A1(n15561), .A2(n15540), .ZN(n7872) );
  INV_X1 U8050 ( .A(n12310), .ZN(n8219) );
  AND2_X1 U8051 ( .A1(n13323), .A2(n11593), .ZN(n8236) );
  NAND2_X1 U8052 ( .A1(n7863), .A2(n7862), .ZN(n11203) );
  NAND2_X1 U8053 ( .A1(n7857), .A2(n7856), .ZN(n13021) );
  NAND2_X1 U8054 ( .A1(n13021), .A2(n13022), .ZN(n10875) );
  OR2_X1 U8055 ( .A1(n12983), .A2(n13341), .ZN(n10870) );
  INV_X1 U8056 ( .A(n13027), .ZN(n13028) );
  NAND2_X1 U8057 ( .A1(n7597), .A2(n7596), .ZN(n15803) );
  INV_X1 U8058 ( .A(n7919), .ZN(n7918) );
  NAND2_X1 U8059 ( .A1(n8485), .A2(n7920), .ZN(n7921) );
  AND2_X1 U8060 ( .A1(n10115), .A2(n14606), .ZN(n8106) );
  OR2_X1 U8061 ( .A1(n8484), .A2(n14425), .ZN(n8487) );
  NAND2_X1 U8062 ( .A1(n8485), .A2(n8486), .ZN(n8257) );
  AND2_X1 U8063 ( .A1(n7942), .A2(SI_16_), .ZN(n7940) );
  INV_X1 U8064 ( .A(n8476), .ZN(n8277) );
  NAND2_X1 U8065 ( .A1(n8475), .A2(SI_13_), .ZN(n8476) );
  OAI21_X1 U8066 ( .B1(n8713), .B2(n8730), .A(n7791), .ZN(n8750) );
  INV_X1 U8067 ( .A(n8250), .ZN(n8249) );
  OAI21_X1 U8068 ( .B1(n8671), .B2(n8251), .A(n8456), .ZN(n8250) );
  INV_X1 U8069 ( .A(n8452), .ZN(n8251) );
  NAND2_X1 U8070 ( .A1(n7634), .A2(n7633), .ZN(n8435) );
  OR2_X1 U8071 ( .A1(n7778), .A2(n10146), .ZN(n7634) );
  INV_X1 U8072 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n16174) );
  OAI21_X1 U8073 ( .B1(n16226), .B2(n16225), .A(n16224), .ZN(n16229) );
  AND2_X1 U8074 ( .A1(n12550), .A2(n12547), .ZN(n12548) );
  INV_X1 U8075 ( .A(n11499), .ZN(n13425) );
  OR2_X1 U8076 ( .A1(n13536), .A2(n7481), .ZN(n8377) );
  NOR2_X1 U8077 ( .A1(n13536), .A2(n8375), .ZN(n8374) );
  INV_X1 U8078 ( .A(n13490), .ZN(n8375) );
  AND2_X1 U8079 ( .A1(n13498), .A2(n7707), .ZN(n7706) );
  NAND2_X1 U8080 ( .A1(n7711), .A2(n13497), .ZN(n7707) );
  NAND2_X1 U8081 ( .A1(n8361), .A2(n13934), .ZN(n8358) );
  NAND2_X1 U8082 ( .A1(n7727), .A2(n7726), .ZN(n11709) );
  AND2_X1 U8083 ( .A1(n8332), .A2(n11505), .ZN(n7726) );
  NAND2_X1 U8084 ( .A1(n7720), .A2(n7718), .ZN(n12549) );
  XNOR2_X1 U8085 ( .A(n11499), .B(n12798), .ZN(n11500) );
  NAND2_X1 U8086 ( .A1(n7724), .A2(n7723), .ZN(n7725) );
  INV_X1 U8087 ( .A(n11195), .ZN(n7723) );
  INV_X1 U8088 ( .A(n11196), .ZN(n7724) );
  AOI21_X1 U8089 ( .B1(n13460), .B2(n13382), .A(n13934), .ZN(n13583) );
  NAND2_X1 U8090 ( .A1(n7730), .A2(n10957), .ZN(n11232) );
  NAND2_X1 U8091 ( .A1(n10977), .A2(n7898), .ZN(n7730) );
  OR2_X1 U8092 ( .A1(n11231), .A2(n7908), .ZN(n7907) );
  OR2_X1 U8093 ( .A1(n11232), .A2(n7908), .ZN(n7904) );
  NAND2_X1 U8094 ( .A1(n11232), .A2(n7906), .ZN(n7901) );
  AND2_X1 U8095 ( .A1(n11231), .A2(n7908), .ZN(n7906) );
  NOR2_X1 U8096 ( .A1(n11766), .A2(n11765), .ZN(n11886) );
  OR2_X1 U8097 ( .A1(n11767), .A2(n16586), .ZN(n7900) );
  NAND2_X1 U8098 ( .A1(n12493), .A2(n12494), .ZN(n13631) );
  OR2_X1 U8099 ( .A1(n13614), .A2(n13613), .ZN(n7912) );
  NAND2_X1 U8100 ( .A1(n7912), .A2(n7911), .ZN(n7910) );
  NAND2_X1 U8101 ( .A1(n13649), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7911) );
  NOR2_X1 U8102 ( .A1(n13651), .A2(n13650), .ZN(n13683) );
  NAND2_X1 U8103 ( .A1(n9572), .A2(n14505), .ZN(n9967) );
  INV_X1 U8104 ( .A(n9952), .ZN(n9572) );
  AOI21_X1 U8105 ( .B1(n7992), .B2(n7996), .A(n7991), .ZN(n7990) );
  NOR2_X1 U8106 ( .A1(n13801), .A2(n13602), .ZN(n7991) );
  NAND2_X1 U8107 ( .A1(n13818), .A2(n13817), .ZN(n7986) );
  AND2_X1 U8108 ( .A1(n12874), .A2(n12871), .ZN(n13864) );
  NOR2_X1 U8109 ( .A1(n13875), .A2(n13876), .ZN(n10019) );
  INV_X1 U8110 ( .A(n13884), .ZN(n14031) );
  AOI21_X1 U8111 ( .B1(n7977), .B2(n7979), .A(n7976), .ZN(n7975) );
  INV_X1 U8112 ( .A(n12820), .ZN(n7976) );
  CLKBUF_X1 U8113 ( .A(n12240), .Z(n7607) );
  AND4_X1 U8114 ( .A1(n9710), .A2(n9709), .A3(n9708), .A4(n9707), .ZN(n12544)
         );
  INV_X1 U8115 ( .A(n13967), .ZN(n13880) );
  NAND2_X1 U8116 ( .A1(n10045), .A2(n12910), .ZN(n13970) );
  INV_X1 U8117 ( .A(n10000), .ZN(n12924) );
  INV_X1 U8118 ( .A(n13878), .ZN(n13973) );
  NAND2_X1 U8119 ( .A1(n10050), .A2(n9479), .ZN(n14052) );
  INV_X1 U8120 ( .A(n13970), .ZN(n13954) );
  NAND2_X1 U8121 ( .A1(n7519), .A2(n7603), .ZN(n16444) );
  INV_X1 U8122 ( .A(n9626), .ZN(n7603) );
  NAND2_X1 U8123 ( .A1(n10059), .A2(n10079), .ZN(n10237) );
  NAND2_X1 U8124 ( .A1(n9555), .A2(n8381), .ZN(n9575) );
  AND2_X1 U8125 ( .A1(n8345), .A2(n7622), .ZN(n7621) );
  AND2_X1 U8126 ( .A1(n7988), .A2(n9556), .ZN(n7622) );
  NAND2_X1 U8127 ( .A1(n9949), .A2(n9542), .ZN(n9962) );
  INV_X1 U8128 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7987) );
  AOI21_X1 U8129 ( .B1(n8151), .B2(n15132), .A(n9933), .ZN(n8148) );
  NAND2_X1 U8130 ( .A1(n8171), .A2(n8169), .ZN(n9906) );
  AOI21_X1 U8131 ( .B1(n7559), .B2(n9882), .A(n8170), .ZN(n8169) );
  INV_X1 U8132 ( .A(n9528), .ZN(n8170) );
  OR2_X1 U8133 ( .A1(n9881), .A2(n9882), .ZN(n8172) );
  NAND2_X1 U8134 ( .A1(n9470), .A2(n9548), .ZN(n9473) );
  NAND2_X1 U8135 ( .A1(n9822), .A2(n8158), .ZN(n8157) );
  NOR2_X1 U8136 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n10389), .ZN(n8166) );
  INV_X1 U8137 ( .A(n8163), .ZN(n8162) );
  OAI21_X1 U8138 ( .B1(n7460), .B2(n10492), .A(n8164), .ZN(n8163) );
  NAND2_X1 U8139 ( .A1(n9762), .A2(n7460), .ZN(n8168) );
  NAND2_X1 U8140 ( .A1(n9762), .A2(n9514), .ZN(n8161) );
  NAND2_X1 U8141 ( .A1(n9728), .A2(n9509), .ZN(n9744) );
  INV_X1 U8142 ( .A(n9698), .ZN(n9503) );
  INV_X1 U8143 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9504) );
  NAND2_X1 U8144 ( .A1(n9684), .A2(n9502), .ZN(n9699) );
  NAND2_X1 U8145 ( .A1(n9500), .A2(n9499), .ZN(n9682) );
  AND2_X1 U8146 ( .A1(n9492), .A2(n9491), .ZN(n9637) );
  NOR2_X1 U8147 ( .A1(n11047), .A2(n8048), .ZN(n8047) );
  NAND2_X1 U8148 ( .A1(n10723), .A2(n8649), .ZN(n8666) );
  INV_X1 U8149 ( .A(n8927), .ZN(n8039) );
  NOR2_X1 U8150 ( .A1(n14687), .A2(n8043), .ZN(n8042) );
  INV_X1 U8151 ( .A(n8901), .ZN(n8043) );
  OR2_X1 U8152 ( .A1(n8777), .A2(n10368), .ZN(n8820) );
  OAI21_X2 U8153 ( .B1(n11460), .B2(n8035), .A(n8033), .ZN(n14629) );
  INV_X1 U8154 ( .A(n8036), .ZN(n8035) );
  AOI21_X1 U8155 ( .B1(n8036), .B2(n8034), .A(n7518), .ZN(n8033) );
  NOR2_X1 U8156 ( .A1(n11694), .A2(n8037), .ZN(n8036) );
  NAND2_X1 U8157 ( .A1(n14618), .A2(n8955), .ZN(n8979) );
  NAND2_X1 U8158 ( .A1(n14735), .A2(n14884), .ZN(n8600) );
  AOI21_X1 U8159 ( .B1(n14629), .B2(n14626), .A(n14624), .ZN(n12087) );
  NAND2_X1 U8160 ( .A1(n12132), .A2(n8026), .ZN(n8025) );
  INV_X1 U8161 ( .A(n8828), .ZN(n8026) );
  OR2_X1 U8162 ( .A1(n8620), .A2(n10590), .ZN(n8595) );
  INV_X1 U8163 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n12129) );
  NAND2_X1 U8164 ( .A1(n9312), .A2(n9311), .ZN(n14804) );
  NAND2_X1 U8165 ( .A1(n9323), .A2(n9322), .ZN(n14810) );
  NAND2_X1 U8166 ( .A1(n7592), .A2(n9356), .ZN(n9323) );
  INV_X1 U8167 ( .A(n15975), .ZN(n7592) );
  OR2_X1 U8168 ( .A1(n14837), .A2(n8075), .ZN(n8074) );
  NAND2_X1 U8169 ( .A1(n14822), .A2(n8076), .ZN(n8075) );
  NAND2_X1 U8170 ( .A1(n7427), .A2(n15016), .ZN(n14844) );
  NAND2_X1 U8171 ( .A1(n8056), .A2(n7748), .ZN(n7747) );
  INV_X1 U8172 ( .A(n14891), .ZN(n7748) );
  OR2_X1 U8173 ( .A1(n14881), .A2(n7749), .ZN(n7743) );
  AND2_X1 U8174 ( .A1(n9013), .A2(n9012), .ZN(n14870) );
  AND2_X1 U8175 ( .A1(n9061), .A2(n9060), .ZN(n14871) );
  NOR2_X1 U8176 ( .A1(n14891), .A2(n8130), .ZN(n8129) );
  INV_X1 U8177 ( .A(n12709), .ZN(n8130) );
  NAND2_X1 U8178 ( .A1(n14910), .A2(n12681), .ZN(n14896) );
  OAI21_X1 U8179 ( .B1(n14946), .B2(n12678), .A(n12679), .ZN(n14939) );
  NAND2_X1 U8180 ( .A1(n12704), .A2(n12703), .ZN(n14929) );
  NAND2_X1 U8181 ( .A1(n12641), .A2(n12642), .ZN(n12674) );
  OR2_X1 U8182 ( .A1(n8054), .A2(n8053), .ZN(n8052) );
  INV_X1 U8183 ( .A(n12586), .ZN(n8053) );
  NAND2_X1 U8184 ( .A1(n12568), .A2(n8054), .ZN(n12587) );
  NAND2_X1 U8185 ( .A1(n12072), .A2(n8146), .ZN(n12190) );
  NAND2_X1 U8186 ( .A1(n8066), .A2(n8064), .ZN(n12192) );
  NOR2_X1 U8187 ( .A1(n12073), .A2(n8065), .ZN(n8064) );
  INV_X1 U8188 ( .A(n8067), .ZN(n8065) );
  INV_X1 U8189 ( .A(n14727), .ZN(n12065) );
  INV_X1 U8190 ( .A(n14911), .ZN(n14951) );
  OR2_X1 U8191 ( .A1(n12032), .A2(n12033), .ZN(n12030) );
  OR2_X1 U8192 ( .A1(n8071), .A2(n8070), .ZN(n7772) );
  INV_X1 U8193 ( .A(n11352), .ZN(n8070) );
  XNOR2_X1 U8194 ( .A(n11934), .B(n14730), .ZN(n11918) );
  INV_X1 U8195 ( .A(n14953), .ZN(n14913) );
  AND2_X1 U8196 ( .A1(n10269), .A2(n10311), .ZN(n14911) );
  NAND2_X1 U8197 ( .A1(n9340), .A2(n9339), .ZN(n15005) );
  NAND2_X1 U8198 ( .A1(n9359), .A2(n9358), .ZN(n15011) );
  NAND2_X1 U8199 ( .A1(n8554), .A2(n8553), .ZN(n15057) );
  NAND2_X1 U8200 ( .A1(n8775), .A2(n8774), .ZN(n12223) );
  AND2_X1 U8201 ( .A1(n8539), .A2(n8509), .ZN(n8416) );
  INV_X1 U8202 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8539) );
  NAND2_X1 U8203 ( .A1(n8871), .A2(n7438), .ZN(n8508) );
  NAND2_X1 U8204 ( .A1(n8522), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8529) );
  OR2_X1 U8205 ( .A1(n8654), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n8690) );
  NAND2_X1 U8206 ( .A1(n10119), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10215) );
  INV_X1 U8207 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n10214) );
  AND2_X1 U8208 ( .A1(n7530), .A2(n10891), .ZN(n7697) );
  NAND2_X1 U8209 ( .A1(n11612), .A2(n11611), .ZN(n8115) );
  INV_X1 U8210 ( .A(n8098), .ZN(n8095) );
  AND2_X1 U8211 ( .A1(n15228), .A2(n8099), .ZN(n8098) );
  NAND2_X1 U8212 ( .A1(n15343), .A2(n15341), .ZN(n8099) );
  NAND2_X1 U8213 ( .A1(n11285), .A2(n11284), .ZN(n8105) );
  NAND2_X1 U8214 ( .A1(n15185), .A2(n15186), .ZN(n8113) );
  NAND2_X1 U8215 ( .A1(n10782), .A2(n10781), .ZN(n7699) );
  NAND2_X1 U8216 ( .A1(n15206), .A2(n15205), .ZN(n7696) );
  NAND2_X1 U8217 ( .A1(n8105), .A2(n8103), .ZN(n11415) );
  NOR2_X1 U8218 ( .A1(n11301), .A2(n8104), .ZN(n8103) );
  INV_X1 U8219 ( .A(n11289), .ZN(n8104) );
  NOR2_X1 U8220 ( .A1(n15311), .A2(n8112), .ZN(n8111) );
  INV_X1 U8221 ( .A(n15183), .ZN(n8112) );
  NAND2_X1 U8222 ( .A1(n15242), .A2(n15243), .ZN(n15241) );
  NAND2_X1 U8223 ( .A1(n15319), .A2(n15320), .ZN(n15318) );
  AND2_X1 U8224 ( .A1(n15331), .A2(n8085), .ZN(n8084) );
  NAND2_X1 U8225 ( .A1(n8088), .A2(n8086), .ZN(n8085) );
  INV_X1 U8226 ( .A(n8089), .ZN(n8086) );
  INV_X1 U8227 ( .A(n8088), .ZN(n8087) );
  NOR2_X1 U8228 ( .A1(n8090), .A2(n15294), .ZN(n8089) );
  NOR2_X1 U8229 ( .A1(n15288), .A2(n7439), .ZN(n8090) );
  AOI21_X1 U8230 ( .B1(n8089), .B2(n7439), .A(n7562), .ZN(n8088) );
  NAND3_X1 U8231 ( .A1(n10783), .A2(n7699), .A3(n7568), .ZN(n7698) );
  NAND2_X1 U8232 ( .A1(n15218), .A2(n15217), .ZN(n8101) );
  AND2_X1 U8233 ( .A1(n7688), .A2(n7687), .ZN(n8102) );
  INV_X1 U8234 ( .A(n7690), .ZN(n7687) );
  OAI21_X1 U8235 ( .B1(n13124), .B2(n13128), .A(n12579), .ZN(n15501) );
  NAND2_X1 U8236 ( .A1(n12975), .A2(n12974), .ZN(n15526) );
  OR2_X1 U8237 ( .A1(n15975), .A2(n12973), .ZN(n12975) );
  AND2_X1 U8238 ( .A1(n7808), .A2(n7806), .ZN(n7812) );
  NAND2_X1 U8239 ( .A1(n7820), .A2(n7807), .ZN(n7806) );
  NAND2_X1 U8240 ( .A1(n7817), .A2(n7813), .ZN(n7808) );
  INV_X1 U8241 ( .A(n15624), .ZN(n7807) );
  NAND2_X1 U8242 ( .A1(n7817), .A2(n7820), .ZN(n7815) );
  OAI211_X1 U8243 ( .C1(n7445), .C2(n7781), .A(n7779), .B(n7938), .ZN(n7937)
         );
  NAND2_X1 U8244 ( .A1(n15578), .A2(n15577), .ZN(n7938) );
  NOR2_X1 U8245 ( .A1(n7880), .A2(n15664), .ZN(n7876) );
  OR2_X1 U8246 ( .A1(n15575), .A2(n8233), .ZN(n8228) );
  INV_X1 U8247 ( .A(n15574), .ZN(n8233) );
  INV_X1 U8248 ( .A(n15575), .ZN(n15696) );
  INV_X1 U8249 ( .A(n15725), .ZN(n7874) );
  NAND2_X1 U8250 ( .A1(n15713), .A2(n15726), .ZN(n15716) );
  INV_X1 U8251 ( .A(n15733), .ZN(n7774) );
  NAND2_X1 U8252 ( .A1(n13157), .A2(n13156), .ZN(n15746) );
  NAND2_X1 U8253 ( .A1(n13137), .A2(n13136), .ZN(n15778) );
  OAI21_X1 U8254 ( .B1(n15541), .B2(n15559), .A(n7872), .ZN(n15817) );
  NAND2_X1 U8255 ( .A1(n15817), .A2(n15816), .ZN(n15815) );
  NAND2_X1 U8256 ( .A1(n12020), .A2(n12019), .ZN(n12021) );
  NAND2_X1 U8257 ( .A1(n12004), .A2(n12003), .ZN(n12311) );
  AND2_X1 U8258 ( .A1(n13322), .A2(n11582), .ZN(n7881) );
  INV_X1 U8259 ( .A(n13322), .ZN(n11810) );
  NAND2_X1 U8260 ( .A1(n11055), .A2(n13311), .ZN(n11057) );
  INV_X1 U8261 ( .A(n11174), .ZN(n8206) );
  OAI22_X1 U8262 ( .A1(n7428), .A2(n10469), .B1(n13204), .B2(n10471), .ZN(
        n8178) );
  AND3_X1 U8263 ( .A1(n15607), .A2(n15910), .A3(n15606), .ZN(n15836) );
  NAND2_X1 U8264 ( .A1(n13185), .A2(n13184), .ZN(n15883) );
  NAND2_X1 U8265 ( .A1(n12002), .A2(n12001), .ZN(n15940) );
  NAND2_X1 U8266 ( .A1(n11865), .A2(n11864), .ZN(n13086) );
  OAI22_X1 U8267 ( .A1(n10392), .A2(P1_D_REG_0__SCAN_IN), .B1(n10391), .B2(
        n10390), .ZN(n11053) );
  AOI21_X1 U8268 ( .B1(n9338), .B2(n9337), .A(n9304), .ZN(n9316) );
  XNOR2_X1 U8269 ( .A(n9355), .B(n9354), .ZN(n13371) );
  INV_X1 U8270 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n10220) );
  NAND2_X1 U8271 ( .A1(n8260), .A2(n9069), .ZN(n9295) );
  NAND2_X1 U8272 ( .A1(n9048), .A2(n8264), .ZN(n8260) );
  NOR2_X1 U8273 ( .A1(n10132), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n10134) );
  NAND2_X1 U8274 ( .A1(n13203), .A2(n8960), .ZN(n8983) );
  XNOR2_X1 U8275 ( .A(n8981), .B(n14417), .ZN(n13203) );
  NAND2_X1 U8276 ( .A1(n8672), .A2(n8671), .ZN(n8674) );
  AND2_X1 U8277 ( .A1(n8652), .A2(n7915), .ZN(n10784) );
  AND2_X1 U8278 ( .A1(n7738), .A2(n7740), .ZN(n7915) );
  AND2_X1 U8279 ( .A1(n8611), .A2(n8569), .ZN(n10494) );
  NOR2_X1 U8280 ( .A1(n16354), .A2(n16355), .ZN(n16222) );
  AOI21_X1 U8281 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n16288), .A(n16287), .ZN(
        n16301) );
  NOR2_X1 U8282 ( .A1(n16286), .A2(n16285), .ZN(n16287) );
  NAND2_X1 U8283 ( .A1(n9919), .A2(n9918), .ZN(n13811) );
  AND4_X1 U8284 ( .A1(n9743), .A2(n9742), .A3(n9741), .A4(n9740), .ZN(n13971)
         );
  NAND2_X1 U8285 ( .A1(n12549), .A2(n12548), .ZN(n12616) );
  INV_X1 U8286 ( .A(n13892), .ZN(n13868) );
  NAND2_X1 U8287 ( .A1(n9874), .A2(n9873), .ZN(n14027) );
  OR2_X1 U8288 ( .A1(n12389), .A2(n12388), .ZN(n12390) );
  NOR2_X1 U8289 ( .A1(n11035), .A2(n11036), .ZN(n11193) );
  NAND2_X1 U8290 ( .A1(n9898), .A2(n9897), .ZN(n14020) );
  INV_X1 U8291 ( .A(n13912), .ZN(n14039) );
  NAND2_X1 U8292 ( .A1(n9845), .A2(n9844), .ZN(n13896) );
  INV_X1 U8293 ( .A(n14123), .ZN(n13597) );
  NAND2_X1 U8294 ( .A1(n10733), .A2(n10732), .ZN(n13599) );
  AOI21_X1 U8295 ( .B1(n12958), .B2(n12765), .A(n7514), .ZN(n8174) );
  INV_X1 U8296 ( .A(n12544), .ZN(n13603) );
  INV_X1 U8297 ( .A(n12388), .ZN(n12394) );
  NAND2_X1 U8298 ( .A1(n7909), .A2(n7493), .ZN(n7737) );
  INV_X1 U8299 ( .A(n7640), .ZN(n13617) );
  AND2_X1 U8300 ( .A1(n9780), .A2(n9779), .ZN(n13961) );
  INV_X1 U8301 ( .A(n13940), .ZN(n13981) );
  AND3_X1 U8302 ( .A1(n9771), .A2(n9770), .A3(n9769), .ZN(n14060) );
  NAND2_X1 U8303 ( .A1(n12135), .A2(n8828), .ZN(n8023) );
  AND2_X1 U8304 ( .A1(n10661), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14700) );
  NAND2_X1 U8305 ( .A1(n8875), .A2(n8874), .ZN(n15073) );
  AND2_X1 U8306 ( .A1(n14662), .A2(n8929), .ZN(n8030) );
  NAND2_X1 U8307 ( .A1(n12087), .A2(n8826), .ZN(n12135) );
  XNOR2_X1 U8308 ( .A(n8979), .B(n8977), .ZN(n14672) );
  NAND2_X1 U8309 ( .A1(n8912), .A2(n8911), .ZN(n15062) );
  AND2_X1 U8310 ( .A1(n9039), .A2(n9038), .ZN(n14695) );
  NAND2_X1 U8311 ( .A1(n8854), .A2(n8853), .ZN(n15078) );
  OR2_X1 U8312 ( .A1(n9442), .A2(n9407), .ZN(n9413) );
  NAND2_X1 U8313 ( .A1(n9085), .A2(n9084), .ZN(n14861) );
  INV_X1 U8314 ( .A(n14871), .ZN(n14838) );
  INV_X1 U8315 ( .A(n14695), .ZN(n14860) );
  INV_X1 U8316 ( .A(n14870), .ZN(n14714) );
  NAND4_X1 U8317 ( .A1(n8624), .A2(n8623), .A3(n8622), .A4(n8621), .ZN(n14733)
         );
  OR2_X1 U8318 ( .A1(n8620), .A2(n10285), .ZN(n8623) );
  NAND2_X1 U8319 ( .A1(n8805), .A2(n8804), .ZN(n16606) );
  AND2_X1 U8320 ( .A1(n10449), .A2(n12727), .ZN(n16507) );
  OR2_X1 U8321 ( .A1(n16522), .A2(n11786), .ZN(n16515) );
  AND2_X1 U8322 ( .A1(n16040), .A2(n9131), .ZN(n16511) );
  INV_X1 U8323 ( .A(n14954), .ZN(n16522) );
  NAND2_X1 U8324 ( .A1(n10391), .A2(n10139), .ZN(n10410) );
  INV_X1 U8325 ( .A(n15614), .ZN(n15653) );
  NAND2_X1 U8326 ( .A1(n12315), .A2(n12314), .ZN(n13102) );
  NAND2_X1 U8327 ( .A1(n13221), .A2(n13220), .ZN(n15867) );
  AND4_X1 U8328 ( .A1(n10509), .A2(n10508), .A3(n10507), .A4(n10506), .ZN(
        n10876) );
  INV_X1 U8329 ( .A(n15778), .ZN(n15905) );
  NAND2_X1 U8330 ( .A1(n13265), .A2(n13264), .ZN(n15847) );
  OAI21_X1 U8331 ( .B1(n13365), .B2(n7463), .A(n7661), .ZN(n7660) );
  INV_X1 U8332 ( .A(n7662), .ZN(n7661) );
  NAND2_X1 U8333 ( .A1(n8190), .A2(n8188), .ZN(n15888) );
  NOR2_X1 U8334 ( .A1(n15741), .A2(n8189), .ZN(n8188) );
  INV_X1 U8335 ( .A(n15548), .ZN(n8189) );
  NAND2_X1 U8336 ( .A1(n13131), .A2(n13130), .ZN(n15909) );
  NAND2_X1 U8337 ( .A1(n8226), .A2(n11567), .ZN(n11569) );
  NAND2_X1 U8338 ( .A1(n15582), .A2(n8200), .ZN(n8199) );
  INV_X1 U8339 ( .A(n15582), .ZN(n8201) );
  NAND2_X1 U8340 ( .A1(n15827), .A2(n7936), .ZN(n7935) );
  INV_X1 U8341 ( .A(n15831), .ZN(n7936) );
  OR2_X1 U8342 ( .A1(n16570), .A2(n8203), .ZN(n8202) );
  INV_X1 U8343 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8203) );
  OAI211_X1 U8344 ( .C1(n15843), .C2(n16435), .A(n15842), .B(n15841), .ZN(
        n15949) );
  NAND2_X1 U8345 ( .A1(n8326), .A2(n7501), .ZN(n15969) );
  INV_X1 U8346 ( .A(n8329), .ZN(n8327) );
  INV_X1 U8347 ( .A(n12983), .ZN(n15997) );
  NOR2_X1 U8348 ( .A1(n16254), .A2(n16253), .ZN(n16255) );
  OAI21_X1 U8349 ( .B1(n16304), .B2(n16305), .A(n7893), .ZN(n7892) );
  INV_X1 U8350 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7893) );
  NOR2_X1 U8351 ( .A1(n16317), .A2(n16316), .ZN(n16318) );
  NAND2_X1 U8352 ( .A1(n16347), .A2(n16346), .ZN(n16348) );
  OAI21_X1 U8353 ( .B1(n16347), .B2(n16346), .A(n7887), .ZN(n7886) );
  INV_X1 U8354 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n7887) );
  NAND2_X1 U8355 ( .A1(n8288), .A2(n13079), .ZN(n8292) );
  NAND2_X1 U8356 ( .A1(n8289), .A2(n13080), .ZN(n8288) );
  NAND2_X1 U8357 ( .A1(n8292), .A2(n8287), .ZN(n8286) );
  NAND2_X1 U8358 ( .A1(n13081), .A2(n13076), .ZN(n8287) );
  NAND2_X1 U8359 ( .A1(n8293), .A2(n13081), .ZN(n8290) );
  INV_X1 U8360 ( .A(n8292), .ZN(n8293) );
  INV_X1 U8361 ( .A(n9171), .ZN(n7594) );
  NAND2_X1 U8362 ( .A1(n8295), .A2(n8294), .ZN(n13093) );
  NAND2_X1 U8363 ( .A1(n13087), .A2(n13089), .ZN(n8294) );
  NOR2_X1 U8364 ( .A1(n9195), .A2(n9193), .ZN(n7854) );
  NAND2_X1 U8365 ( .A1(n8301), .A2(n8300), .ZN(n13115) );
  NAND2_X1 U8366 ( .A1(n13106), .A2(n13108), .ZN(n8300) );
  AND2_X1 U8367 ( .A1(n9208), .A2(n8386), .ZN(n8385) );
  NAND2_X1 U8368 ( .A1(n8304), .A2(n8303), .ZN(n13147) );
  NAND2_X1 U8369 ( .A1(n13132), .A2(n13134), .ZN(n8303) );
  NAND2_X1 U8370 ( .A1(n8409), .A2(n8408), .ZN(n8407) );
  INV_X1 U8371 ( .A(n9233), .ZN(n8408) );
  INV_X1 U8372 ( .A(n9234), .ZN(n8409) );
  NAND2_X1 U8373 ( .A1(n13165), .A2(n8320), .ZN(n8319) );
  OAI21_X1 U8374 ( .B1(n9230), .B2(n9229), .A(n9228), .ZN(n9235) );
  OAI21_X1 U8375 ( .B1(n9221), .B2(n8391), .A(n8389), .ZN(n9230) );
  OAI21_X1 U8376 ( .B1(n9221), .B2(n8394), .A(n7510), .ZN(n9228) );
  NOR2_X1 U8377 ( .A1(n7614), .A2(n9241), .ZN(n7613) );
  INV_X1 U8378 ( .A(n8407), .ZN(n7614) );
  AND2_X1 U8379 ( .A1(n9233), .A2(n9234), .ZN(n8410) );
  INV_X1 U8380 ( .A(n9249), .ZN(n7840) );
  AND2_X1 U8381 ( .A1(n9242), .A2(n8418), .ZN(n7586) );
  NAND2_X1 U8382 ( .A1(n8419), .A2(n9245), .ZN(n8418) );
  OAI21_X1 U8383 ( .B1(n9235), .B2(n8410), .A(n7613), .ZN(n9242) );
  INV_X1 U8384 ( .A(n7521), .ZN(n8419) );
  INV_X1 U8385 ( .A(n7552), .ZN(n8412) );
  NOR2_X1 U8386 ( .A1(n9250), .A2(n7840), .ZN(n7838) );
  AND2_X1 U8387 ( .A1(n9250), .A2(n7840), .ZN(n7839) );
  NAND2_X1 U8388 ( .A1(n13180), .A2(n7681), .ZN(n7682) );
  NAND2_X1 U8389 ( .A1(n13193), .A2(n13195), .ZN(n8307) );
  OAI22_X1 U8390 ( .A1(n13206), .A2(n7654), .B1(n13207), .B2(n7653), .ZN(
        n13224) );
  INV_X1 U8391 ( .A(n13205), .ZN(n7653) );
  NOR2_X1 U8392 ( .A1(n13208), .A2(n13205), .ZN(n7654) );
  NAND2_X1 U8393 ( .A1(n8308), .A2(n8307), .ZN(n13206) );
  NAND2_X1 U8394 ( .A1(n7552), .A2(n8414), .ZN(n8413) );
  NAND2_X1 U8395 ( .A1(n9258), .A2(n9257), .ZN(n7590) );
  NAND2_X1 U8396 ( .A1(n13224), .A2(n13225), .ZN(n13223) );
  NAND2_X1 U8397 ( .A1(n7587), .A2(n7588), .ZN(n9265) );
  OR2_X1 U8398 ( .A1(n9258), .A2(n9257), .ZN(n7587) );
  NAND2_X1 U8399 ( .A1(n7590), .A2(n7589), .ZN(n7588) );
  INV_X1 U8400 ( .A(n9256), .ZN(n7589) );
  INV_X1 U8401 ( .A(n9263), .ZN(n7830) );
  INV_X1 U8402 ( .A(n9268), .ZN(n8422) );
  INV_X1 U8403 ( .A(n9269), .ZN(n8423) );
  OAI21_X1 U8404 ( .B1(n7829), .B2(n7828), .A(n8421), .ZN(n9274) );
  NAND2_X1 U8405 ( .A1(n8423), .A2(n8422), .ZN(n8421) );
  AOI21_X1 U8406 ( .B1(n9265), .B2(n9264), .A(n7830), .ZN(n7829) );
  OAI21_X1 U8407 ( .B1(n9265), .B2(n9264), .A(n7513), .ZN(n7828) );
  NAND2_X1 U8408 ( .A1(n8312), .A2(n8311), .ZN(n13268) );
  NAND2_X1 U8409 ( .A1(n13253), .A2(n13255), .ZN(n8311) );
  INV_X1 U8410 ( .A(n13293), .ZN(n8323) );
  NAND2_X1 U8411 ( .A1(n7523), .A2(n7454), .ZN(n7673) );
  AND2_X1 U8412 ( .A1(n13876), .A2(n13887), .ZN(n12942) );
  NOR2_X1 U8413 ( .A1(n12934), .A2(n8008), .ZN(n8005) );
  INV_X1 U8414 ( .A(n10008), .ZN(n8008) );
  NAND2_X1 U8415 ( .A1(n10008), .A2(n8007), .ZN(n8006) );
  INV_X1 U8416 ( .A(n10007), .ZN(n8007) );
  OR2_X1 U8417 ( .A1(n10237), .A2(P3_D_REG_0__SCAN_IN), .ZN(n11028) );
  NAND2_X1 U8418 ( .A1(n9283), .A2(n9284), .ZN(n8399) );
  NAND2_X1 U8419 ( .A1(n8402), .A2(n8401), .ZN(n8400) );
  INV_X1 U8420 ( .A(n9284), .ZN(n8402) );
  NOR2_X1 U8421 ( .A1(n7548), .A2(n8397), .ZN(n8396) );
  INV_X1 U8422 ( .A(n8399), .ZN(n8397) );
  INV_X1 U8423 ( .A(n14726), .ZN(n8069) );
  OR2_X1 U8424 ( .A1(n15876), .A2(n15554), .ZN(n15576) );
  INV_X1 U8425 ( .A(n8262), .ZN(n8261) );
  OAI21_X1 U8426 ( .B1(n8264), .B2(n8263), .A(n9294), .ZN(n8262) );
  INV_X1 U8427 ( .A(n9069), .ZN(n8263) );
  NOR2_X1 U8428 ( .A1(n7922), .A2(n8902), .ZN(n7920) );
  OAI21_X1 U8429 ( .B1(n7922), .B2(n7927), .A(n8281), .ZN(n7919) );
  AOI21_X1 U8430 ( .B1(n8283), .B2(n8282), .A(n7553), .ZN(n8281) );
  INV_X1 U8431 ( .A(n8938), .ZN(n8282) );
  INV_X1 U8432 ( .A(n8934), .ZN(n8937) );
  INV_X1 U8433 ( .A(n8551), .ZN(n7927) );
  AND2_X1 U8434 ( .A1(n8482), .A2(n7801), .ZN(n7800) );
  INV_X1 U8435 ( .A(n8887), .ZN(n7801) );
  OR2_X1 U8436 ( .A1(n7799), .A2(n8867), .ZN(n7798) );
  INV_X1 U8437 ( .A(n7930), .ZN(n7929) );
  INV_X1 U8438 ( .A(n7791), .ZN(n7790) );
  NOR2_X1 U8439 ( .A1(n8769), .A2(n7931), .ZN(n7930) );
  INV_X1 U8440 ( .A(n8468), .ZN(n7931) );
  NAND2_X1 U8441 ( .A1(n7789), .A2(n8730), .ZN(n7788) );
  OR2_X1 U8442 ( .A1(n8614), .A2(n8444), .ZN(n7742) );
  INV_X1 U8443 ( .A(n8631), .ZN(n8442) );
  NAND2_X1 U8444 ( .A1(n7896), .A2(n7898), .ZN(n10975) );
  NAND2_X1 U8445 ( .A1(n11667), .A2(n11666), .ZN(n7733) );
  NAND2_X1 U8446 ( .A1(n7733), .A2(n11720), .ZN(n11668) );
  NAND2_X1 U8447 ( .A1(n12438), .A2(n12442), .ZN(n12492) );
  NAND2_X1 U8448 ( .A1(n13619), .A2(n13618), .ZN(n7639) );
  NOR2_X1 U8449 ( .A1(n13667), .A2(n7641), .ZN(n13670) );
  NOR2_X1 U8450 ( .A1(n7643), .A2(n7642), .ZN(n7641) );
  INV_X1 U8451 ( .A(n13669), .ZN(n7643) );
  NOR2_X1 U8452 ( .A1(n7995), .A2(n10028), .ZN(n7994) );
  INV_X1 U8453 ( .A(n7996), .ZN(n7995) );
  NOR2_X1 U8454 ( .A1(n10028), .A2(n7999), .ZN(n7992) );
  NAND2_X1 U8455 ( .A1(n9569), .A2(n14497), .ZN(n9920) );
  INV_X1 U8456 ( .A(n9911), .ZN(n9569) );
  OR2_X1 U8457 ( .A1(n9899), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9911) );
  INV_X1 U8458 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n14493) );
  NAND2_X1 U8459 ( .A1(n9563), .A2(n14272), .ZN(n9736) );
  INV_X1 U8460 ( .A(n9722), .ZN(n9563) );
  NAND2_X1 U8461 ( .A1(n13607), .A2(n16444), .ZN(n12800) );
  INV_X1 U8462 ( .A(n11194), .ZN(n7958) );
  INV_X1 U8463 ( .A(n12936), .ZN(n7960) );
  INV_X1 U8464 ( .A(n7978), .ZN(n7977) );
  OAI21_X1 U8465 ( .B1(n12812), .B2(n7979), .A(n12924), .ZN(n7978) );
  INV_X1 U8466 ( .A(n12816), .ZN(n7979) );
  CLKBUF_X1 U8467 ( .A(n11749), .Z(n11947) );
  NAND2_X1 U8468 ( .A1(n12792), .A2(n12927), .ZN(n11626) );
  NOR2_X1 U8469 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), .ZN(
        n7988) );
  AND2_X1 U8470 ( .A1(n9464), .A2(n7729), .ZN(n9807) );
  INV_X1 U8471 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7729) );
  NAND2_X1 U8472 ( .A1(n8165), .A2(n10389), .ZN(n8164) );
  INV_X1 U8473 ( .A(n9514), .ZN(n8165) );
  NAND2_X1 U8474 ( .A1(n10227), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9507) );
  AND2_X1 U8475 ( .A1(n8366), .A2(n8364), .ZN(n9686) );
  NAND2_X1 U8476 ( .A1(n10175), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9496) );
  NAND2_X1 U8477 ( .A1(n10160), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9492) );
  INV_X1 U8478 ( .A(n9624), .ZN(n8366) );
  INV_X1 U8479 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n9455) );
  NAND2_X1 U8480 ( .A1(n9455), .A2(n8368), .ZN(n8367) );
  INV_X1 U8481 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8368) );
  INV_X1 U8482 ( .A(n8768), .ZN(n8037) );
  INV_X1 U8483 ( .A(n11461), .ZN(n8034) );
  NAND2_X1 U8484 ( .A1(n7746), .A2(n7744), .ZN(n14835) );
  AOI21_X1 U8485 ( .B1(n7440), .B2(n7749), .A(n7745), .ZN(n7744) );
  INV_X1 U8486 ( .A(n12689), .ZN(n7745) );
  NAND2_X1 U8487 ( .A1(n7950), .A2(n14877), .ZN(n7949) );
  INV_X1 U8488 ( .A(n7951), .ZN(n7950) );
  NAND2_X1 U8489 ( .A1(n14889), .A2(n7952), .ZN(n7951) );
  NOR2_X1 U8490 ( .A1(n14989), .A2(n15057), .ZN(n12718) );
  NAND2_X1 U8491 ( .A1(n8536), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8892) );
  INV_X1 U8492 ( .A(n8877), .ZN(n8536) );
  AND2_X1 U8493 ( .A1(n7956), .A2(n7955), .ZN(n7954) );
  INV_X1 U8494 ( .A(n12189), .ZN(n8145) );
  NOR2_X1 U8495 ( .A1(n16606), .A2(n12223), .ZN(n7956) );
  NAND2_X1 U8496 ( .A1(n12192), .A2(n12191), .ZN(n12193) );
  AND2_X1 U8497 ( .A1(n12147), .A2(n16573), .ZN(n12078) );
  INV_X1 U8498 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8718) );
  NOR2_X1 U8499 ( .A1(n11923), .A2(n8072), .ZN(n8071) );
  INV_X1 U8500 ( .A(n11348), .ZN(n8072) );
  AND2_X1 U8501 ( .A1(n10995), .A2(n10815), .ZN(n8060) );
  INV_X1 U8502 ( .A(n10818), .ZN(n8062) );
  NAND2_X1 U8503 ( .A1(n14985), .A2(n14995), .ZN(n14989) );
  OR2_X1 U8504 ( .A1(n15073), .A2(n12595), .ZN(n12651) );
  AND2_X1 U8505 ( .A1(n11927), .A2(n16499), .ZN(n11928) );
  INV_X1 U8506 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8500) );
  INV_X1 U8507 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8501) );
  NOR2_X1 U8508 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n8516) );
  INV_X1 U8509 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9125) );
  NAND2_X1 U8510 ( .A1(n9103), .A2(n9102), .ZN(n9124) );
  INV_X1 U8511 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9102) );
  INV_X1 U8512 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8831) );
  OR2_X1 U8513 ( .A1(n13027), .A2(n10338), .ZN(n15136) );
  INV_X1 U8514 ( .A(n13362), .ZN(n7665) );
  NOR2_X1 U8515 ( .A1(n7464), .A2(n7814), .ZN(n7813) );
  NOR2_X1 U8516 ( .A1(n15685), .A2(n15859), .ZN(n8214) );
  NAND2_X1 U8517 ( .A1(n8228), .A2(n15576), .ZN(n8227) );
  NOR2_X1 U8518 ( .A1(n15774), .A2(n15746), .ZN(n15527) );
  OR2_X1 U8519 ( .A1(n13082), .A2(n8213), .ZN(n8212) );
  NAND2_X1 U8520 ( .A1(n7599), .A2(n7598), .ZN(n11981) );
  NOR2_X1 U8521 ( .A1(n8212), .A2(n13086), .ZN(n7598) );
  OR2_X1 U8522 ( .A1(n13078), .A2(n16526), .ZN(n8213) );
  AND2_X1 U8523 ( .A1(n7447), .A2(n11591), .ZN(n8223) );
  NAND2_X1 U8524 ( .A1(n7601), .A2(n7600), .ZN(n10862) );
  INV_X1 U8525 ( .A(n15527), .ZN(n15748) );
  NOR2_X1 U8526 ( .A1(n9070), .A2(n8265), .ZN(n8264) );
  INV_X1 U8527 ( .A(n9047), .ZN(n8265) );
  NAND2_X1 U8528 ( .A1(n8254), .A2(n8252), .ZN(n9020) );
  INV_X1 U8529 ( .A(n8253), .ZN(n8252) );
  OAI21_X1 U8530 ( .B1(n8982), .B2(n8996), .A(n8999), .ZN(n8253) );
  NAND2_X1 U8531 ( .A1(n8107), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10216) );
  AND2_X1 U8532 ( .A1(n8110), .A2(n8109), .ZN(n8108) );
  AOI21_X1 U8533 ( .B1(n8811), .B2(n8276), .A(n7515), .ZN(n8274) );
  INV_X1 U8534 ( .A(n10203), .ZN(n10250) );
  OR2_X1 U8535 ( .A1(n10193), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n10203) );
  INV_X1 U8536 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n14583) );
  AND2_X1 U8537 ( .A1(n8449), .A2(n8448), .ZN(n8650) );
  NAND2_X1 U8538 ( .A1(n7751), .A2(SI_3_), .ZN(n8629) );
  NAND2_X1 U8539 ( .A1(n7755), .A2(n7754), .ZN(n7751) );
  OAI211_X1 U8540 ( .C1(n7755), .C2(n7753), .A(n7752), .B(n7509), .ZN(n8608)
         );
  NOR2_X1 U8541 ( .A1(n7753), .A2(n7671), .ZN(n7750) );
  NAND2_X1 U8542 ( .A1(n7757), .A2(n7756), .ZN(n8568) );
  NAND2_X1 U8543 ( .A1(n7778), .A2(n10493), .ZN(n7756) );
  OR2_X1 U8544 ( .A1(n7778), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7757) );
  INV_X1 U8545 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n16175) );
  INV_X1 U8546 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n16184) );
  NOR2_X1 U8547 ( .A1(n16233), .A2(n16232), .ZN(n16247) );
  NOR2_X1 U8548 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n16231), .ZN(n16232) );
  OAI21_X1 U8549 ( .B1(n16266), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n16265), .ZN(
        n16279) );
  OR2_X1 U8550 ( .A1(n16264), .A2(n16263), .ZN(n16265) );
  OAI21_X1 U8551 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n16282), .A(n16281), .ZN(
        n16286) );
  OR2_X1 U8552 ( .A1(n16280), .A2(n16279), .ZN(n16281) );
  INV_X1 U8553 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n14272) );
  AOI21_X1 U8554 ( .B1(n13453), .B2(n13423), .A(n13427), .ZN(n8341) );
  INV_X1 U8555 ( .A(n8341), .ZN(n8338) );
  AOI21_X1 U8556 ( .B1(n7448), .B2(n8344), .A(n7507), .ZN(n8342) );
  AND2_X1 U8557 ( .A1(n13420), .A2(n13419), .ZN(n13498) );
  NAND2_X1 U8558 ( .A1(n8361), .A2(n13382), .ZN(n8360) );
  NAND2_X1 U8559 ( .A1(n8348), .A2(n8349), .ZN(n13518) );
  AOI22_X1 U8560 ( .A1(n8350), .A2(n8351), .B1(n8352), .B2(n8354), .ZN(n8349)
         );
  INV_X1 U8561 ( .A(n8358), .ZN(n8354) );
  AND2_X1 U8562 ( .A1(n13497), .A2(n13416), .ZN(n13527) );
  INV_X1 U8563 ( .A(n13527), .ZN(n7711) );
  INV_X1 U8564 ( .A(n13795), .ZN(n13531) );
  OAI21_X1 U8565 ( .B1(n13406), .B2(n13405), .A(n13408), .ZN(n13555) );
  AND2_X1 U8566 ( .A1(n13404), .A2(n13403), .ZN(n13554) );
  AND2_X1 U8567 ( .A1(n8376), .A2(n8371), .ZN(n8370) );
  NAND2_X1 U8568 ( .A1(n14140), .A2(n10737), .ZN(n10929) );
  OR2_X1 U8569 ( .A1(n7436), .A2(n10941), .ZN(n9633) );
  OR2_X1 U8570 ( .A1(n7619), .A2(n16428), .ZN(n7735) );
  NAND2_X1 U8571 ( .A1(n7731), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n10977) );
  INV_X1 U8572 ( .A(n10975), .ZN(n7731) );
  OR2_X1 U8573 ( .A1(n9700), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n9715) );
  NAND2_X1 U8574 ( .A1(n7905), .A2(n11385), .ZN(n11403) );
  NAND2_X1 U8575 ( .A1(n11232), .A2(n11231), .ZN(n7905) );
  NOR2_X1 U8576 ( .A1(n7903), .A2(n12280), .ZN(n7902) );
  INV_X1 U8577 ( .A(n7907), .ZN(n7903) );
  NOR2_X1 U8578 ( .A1(n11230), .A2(n7616), .ZN(n7615) );
  INV_X1 U8579 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n7616) );
  NAND2_X1 U8580 ( .A1(n11668), .A2(n7732), .ZN(n11669) );
  OR2_X1 U8581 ( .A1(n7733), .A2(n11720), .ZN(n7732) );
  NOR2_X1 U8582 ( .A1(n11669), .A2(n16542), .ZN(n11726) );
  NAND2_X1 U8583 ( .A1(n11663), .A2(n7635), .ZN(n11721) );
  OR2_X1 U8584 ( .A1(n11665), .A2(n11390), .ZN(n7635) );
  NOR2_X1 U8585 ( .A1(n11726), .A2(n7913), .ZN(n11728) );
  INV_X1 U8586 ( .A(n11668), .ZN(n7913) );
  NAND2_X1 U8587 ( .A1(n7900), .A2(n7488), .ZN(n7899) );
  NAND2_X1 U8588 ( .A1(n11907), .A2(n11908), .ZN(n12438) );
  NAND2_X1 U8589 ( .A1(n7617), .A2(n13628), .ZN(n13630) );
  NAND2_X1 U8590 ( .A1(n13631), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7617) );
  NOR2_X1 U8591 ( .A1(n16369), .A2(n16370), .ZN(n16368) );
  XNOR2_X1 U8592 ( .A(n13610), .B(n13632), .ZN(n16372) );
  AND2_X1 U8593 ( .A1(n13609), .A2(n13608), .ZN(n13610) );
  NOR2_X1 U8594 ( .A1(n13647), .A2(n7644), .ZN(n13667) );
  NAND2_X1 U8595 ( .A1(n7646), .A2(n7645), .ZN(n7644) );
  INV_X1 U8596 ( .A(n13646), .ZN(n7645) );
  INV_X1 U8597 ( .A(n13645), .ZN(n7646) );
  INV_X1 U8598 ( .A(n7910), .ZN(n13660) );
  OR2_X1 U8599 ( .A1(n9967), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9982) );
  NAND2_X1 U8600 ( .A1(n9571), .A2(n9570), .ZN(n9952) );
  INV_X1 U8601 ( .A(n9939), .ZN(n9571) );
  OR2_X1 U8602 ( .A1(n9920), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9928) );
  OR2_X1 U8603 ( .A1(n9928), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9939) );
  NAND2_X1 U8604 ( .A1(n9568), .A2(n14291), .ZN(n9899) );
  INV_X1 U8605 ( .A(n9885), .ZN(n9568) );
  OR2_X1 U8606 ( .A1(n9875), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9885) );
  OR2_X1 U8607 ( .A1(n9846), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9863) );
  NAND2_X1 U8608 ( .A1(n9567), .A2(n14295), .ZN(n9875) );
  INV_X1 U8609 ( .A(n9863), .ZN(n9567) );
  OR2_X1 U8610 ( .A1(n9812), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9832) );
  NAND2_X1 U8611 ( .A1(n9566), .A2(n13511), .ZN(n9846) );
  INV_X1 U8612 ( .A(n9832), .ZN(n9566) );
  AND2_X1 U8613 ( .A1(n12862), .A2(n12860), .ZN(n13907) );
  NAND2_X1 U8614 ( .A1(n10013), .A2(n12848), .ZN(n13933) );
  NAND2_X1 U8615 ( .A1(n9564), .A2(n14493), .ZN(n9796) );
  INV_X1 U8616 ( .A(n9781), .ZN(n9564) );
  NAND2_X1 U8617 ( .A1(n9565), .A2(n14464), .ZN(n9812) );
  INV_X1 U8618 ( .A(n9796), .ZN(n9565) );
  NAND2_X1 U8619 ( .A1(n8011), .A2(n10011), .ZN(n13950) );
  OR2_X1 U8620 ( .A1(n9736), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9752) );
  INV_X1 U8621 ( .A(n7964), .ZN(n7963) );
  NAND2_X1 U8622 ( .A1(n10006), .A2(n12306), .ZN(n12302) );
  OR2_X1 U8623 ( .A1(n9704), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n9722) );
  NAND2_X1 U8624 ( .A1(n9562), .A2(n14273), .ZN(n9704) );
  INV_X1 U8625 ( .A(n9692), .ZN(n9562) );
  OR2_X1 U8626 ( .A1(n9675), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9692) );
  OR2_X1 U8627 ( .A1(n7430), .A2(SI_5_), .ZN(n9661) );
  NAND2_X1 U8628 ( .A1(n11254), .A2(n14472), .ZN(n9663) );
  INV_X1 U8629 ( .A(n12795), .ZN(n12930) );
  NAND2_X1 U8630 ( .A1(n9598), .A2(n11032), .ZN(n11537) );
  NAND2_X1 U8631 ( .A1(n9990), .A2(n12788), .ZN(n12922) );
  CLKBUF_X1 U8632 ( .A(n13748), .Z(n13749) );
  NAND2_X1 U8633 ( .A1(n8009), .A2(n10032), .ZN(n13751) );
  AOI21_X1 U8634 ( .B1(n7984), .B2(n7982), .A(n7981), .ZN(n7980) );
  INV_X1 U8635 ( .A(n7984), .ZN(n7983) );
  INV_X1 U8636 ( .A(n12893), .ZN(n7981) );
  AND2_X1 U8637 ( .A1(n12781), .A2(n12780), .ZN(n13791) );
  OAI21_X1 U8638 ( .B1(n13822), .B2(n7998), .A(n7996), .ZN(n13792) );
  NAND2_X1 U8639 ( .A1(n7986), .A2(n7984), .ZN(n14008) );
  NAND2_X1 U8640 ( .A1(n7967), .A2(n7968), .ZN(n13849) );
  AOI21_X1 U8641 ( .B1(n7971), .B2(n7973), .A(n7969), .ZN(n7968) );
  INV_X1 U8642 ( .A(n12871), .ZN(n7969) );
  AOI21_X1 U8643 ( .B1(n13876), .B2(n8015), .A(n8013), .ZN(n8012) );
  NOR2_X1 U8644 ( .A1(n13871), .A2(n13879), .ZN(n8013) );
  INV_X1 U8645 ( .A(n14052), .ZN(n14015) );
  NAND2_X1 U8646 ( .A1(n13930), .A2(n9787), .ZN(n13949) );
  AND2_X1 U8647 ( .A1(n12844), .A2(n12843), .ZN(n13966) );
  AND4_X1 U8648 ( .A1(n9680), .A2(n9679), .A3(n9678), .A4(n9677), .ZN(n12388)
         );
  NOR2_X1 U8649 ( .A1(n12932), .A2(n8002), .ZN(n8001) );
  INV_X1 U8650 ( .A(n10001), .ZN(n8002) );
  CLKBUF_X1 U8651 ( .A(n12107), .Z(n12108) );
  INV_X1 U8652 ( .A(n12931), .ZN(n12812) );
  NAND2_X1 U8653 ( .A1(n11746), .A2(n12812), .ZN(n11748) );
  INV_X1 U8654 ( .A(n16580), .ZN(n14040) );
  AND2_X1 U8655 ( .A1(n8381), .A2(n8380), .ZN(n8379) );
  INV_X1 U8656 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8380) );
  NOR2_X1 U8657 ( .A1(n9933), .A2(n15132), .ZN(n8150) );
  INV_X1 U8658 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9549) );
  OAI21_X1 U8659 ( .B1(n10074), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n10076) );
  AND2_X1 U8660 ( .A1(n9475), .A2(n10074), .ZN(n12789) );
  AOI21_X1 U8661 ( .B1(n8154), .B2(n8155), .A(n8153), .ZN(n8152) );
  INV_X1 U8662 ( .A(n9523), .ZN(n8153) );
  INV_X1 U8663 ( .A(n8158), .ZN(n8154) );
  INV_X1 U8664 ( .A(n9464), .ZN(n9791) );
  AND2_X1 U8665 ( .A1(n9514), .A2(n9513), .ZN(n9759) );
  AND2_X1 U8666 ( .A1(n9509), .A2(n9508), .ZN(n9729) );
  XNOR2_X1 U8667 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n9698) );
  INV_X1 U8668 ( .A(n9681), .ZN(n7576) );
  NAND2_X1 U8669 ( .A1(n8366), .A2(n9455), .ZN(n9639) );
  AND2_X1 U8670 ( .A1(n9489), .A2(n9488), .ZN(n9622) );
  INV_X1 U8671 ( .A(n8365), .ZN(n9624) );
  XNOR2_X1 U8672 ( .A(n7914), .B(n9616), .ZN(n11097) );
  NAND2_X1 U8673 ( .A1(n7636), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7914) );
  INV_X1 U8674 ( .A(n9615), .ZN(n7636) );
  OR2_X1 U8675 ( .A1(n8697), .A2(n8696), .ZN(n8719) );
  OR2_X1 U8676 ( .A1(n8557), .A2(n14664), .ZN(n8943) );
  INV_X1 U8677 ( .A(n14616), .ZN(n8028) );
  INV_X1 U8678 ( .A(n14654), .ZN(n8020) );
  NAND2_X1 U8679 ( .A1(n8535), .A2(n8534), .ZN(n8837) );
  INV_X1 U8680 ( .A(n8820), .ZN(n8535) );
  NAND2_X1 U8681 ( .A1(n12542), .A2(n8042), .ZN(n14684) );
  NAND2_X1 U8682 ( .A1(n10727), .A2(n8047), .ZN(n11045) );
  AND2_X1 U8683 ( .A1(n8519), .A2(n9405), .ZN(n10269) );
  OR2_X1 U8684 ( .A1(n8858), .A2(n8857), .ZN(n8877) );
  NAND2_X1 U8685 ( .A1(n9376), .A2(n7550), .ZN(n7841) );
  NAND2_X1 U8686 ( .A1(n9376), .A2(n7551), .ZN(n7845) );
  NAND2_X1 U8687 ( .A1(n7851), .A2(n7847), .ZN(n7846) );
  NAND2_X1 U8688 ( .A1(n7850), .A2(n7849), .ZN(n7848) );
  NOR2_X1 U8689 ( .A1(n9389), .A2(n8268), .ZN(n8267) );
  AND2_X1 U8690 ( .A1(n9390), .A2(n9391), .ZN(n8268) );
  NOR2_X1 U8691 ( .A1(n14811), .A2(n14810), .ZN(n14812) );
  NAND2_X1 U8692 ( .A1(n14824), .A2(n12723), .ZN(n14811) );
  AOI21_X1 U8693 ( .B1(n8134), .B2(n8133), .A(n7498), .ZN(n8132) );
  INV_X1 U8694 ( .A(n12714), .ZN(n8133) );
  OAI21_X1 U8695 ( .B1(n14837), .B2(n14821), .A(n8078), .ZN(n8077) );
  XNOR2_X1 U8696 ( .A(n14843), .B(n14861), .ZN(n14834) );
  AND2_X1 U8697 ( .A1(n9078), .A2(n9055), .ZN(n14854) );
  NOR2_X1 U8698 ( .A1(n14918), .A2(n7949), .ZN(n14872) );
  OAI21_X1 U8699 ( .B1(n14899), .B2(n8128), .A(n8126), .ZN(n14866) );
  INV_X1 U8700 ( .A(n8129), .ZN(n8128) );
  AOI21_X1 U8701 ( .B1(n8129), .B2(n8127), .A(n7495), .ZN(n8126) );
  AND2_X1 U8702 ( .A1(n9007), .A2(n9032), .ZN(n14887) );
  NOR2_X1 U8703 ( .A1(n14918), .A2(n15035), .ZN(n14903) );
  NOR2_X1 U8704 ( .A1(n14918), .A2(n7951), .ZN(n14885) );
  NAND2_X1 U8705 ( .A1(n7520), .A2(n7770), .ZN(n14910) );
  INV_X1 U8706 ( .A(n14715), .ZN(n14942) );
  INV_X1 U8707 ( .A(n12718), .ZN(n14969) );
  NAND2_X1 U8708 ( .A1(n7426), .A2(n7583), .ZN(n14968) );
  AOI21_X1 U8709 ( .B1(n7450), .B2(n7762), .A(n7502), .ZN(n7760) );
  NAND2_X1 U8710 ( .A1(n12593), .A2(n7453), .ZN(n12649) );
  OAI21_X1 U8711 ( .B1(n12072), .B2(n8144), .A(n8142), .ZN(n12263) );
  INV_X1 U8712 ( .A(n8143), .ZN(n8142) );
  OAI22_X1 U8713 ( .A1(n8146), .A2(n8144), .B1(n16606), .B2(n14724), .ZN(n8143) );
  OR2_X1 U8714 ( .A1(n12261), .A2(n8145), .ZN(n8144) );
  AND2_X1 U8715 ( .A1(n7765), .A2(n12267), .ZN(n7764) );
  NAND2_X1 U8716 ( .A1(n7766), .A2(n7769), .ZN(n7765) );
  NAND2_X1 U8717 ( .A1(n12078), .A2(n7956), .ZN(n12273) );
  NAND2_X1 U8718 ( .A1(n12078), .A2(n12082), .ZN(n12201) );
  INV_X1 U8719 ( .A(n8140), .ZN(n8139) );
  AOI21_X1 U8720 ( .B1(n8140), .B2(n8138), .A(n7486), .ZN(n8137) );
  AND2_X1 U8721 ( .A1(n8141), .A2(n12069), .ZN(n8140) );
  NOR2_X1 U8722 ( .A1(n12036), .A2(n12095), .ZN(n12147) );
  OR2_X1 U8723 ( .A1(n8719), .A2(n8718), .ZN(n8736) );
  INV_X1 U8724 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8735) );
  OR2_X1 U8725 ( .A1(n8736), .A2(n8735), .ZN(n8756) );
  NAND2_X1 U8726 ( .A1(n7948), .A2(n7947), .ZN(n12036) );
  INV_X1 U8727 ( .A(n14729), .ZN(n12029) );
  NAND2_X1 U8728 ( .A1(n11349), .A2(n8071), .ZN(n11920) );
  NAND2_X1 U8729 ( .A1(n8119), .A2(n8120), .ZN(n11343) );
  AOI21_X1 U8730 ( .B1(n8122), .B2(n8121), .A(n7500), .ZN(n8120) );
  NAND2_X1 U8731 ( .A1(n11349), .A2(n11348), .ZN(n11922) );
  INV_X1 U8732 ( .A(n10610), .ZN(n10604) );
  NAND2_X1 U8733 ( .A1(n8513), .A2(n8512), .ZN(n15053) );
  NAND2_X1 U8734 ( .A1(n8695), .A2(n8694), .ZN(n11548) );
  AND2_X1 U8735 ( .A1(n15121), .A2(n9114), .ZN(n16034) );
  NAND2_X1 U8736 ( .A1(n9105), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9108) );
  INV_X1 U8737 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9107) );
  NAND2_X1 U8738 ( .A1(n9108), .A2(n9107), .ZN(n9110) );
  NAND2_X1 U8739 ( .A1(n9104), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9112) );
  OR2_X1 U8740 ( .A1(n9124), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n9104) );
  INV_X1 U8741 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9111) );
  INV_X1 U8742 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8528) );
  OR2_X1 U8743 ( .A1(n8714), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8732) );
  CLKBUF_X1 U8744 ( .A(n8633), .Z(n8634) );
  INV_X1 U8745 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8492) );
  NOR2_X1 U8746 ( .A1(n12008), .A2(n12007), .ZN(n12321) );
  NAND2_X1 U8747 ( .A1(n12516), .A2(n7497), .ZN(n15148) );
  AOI21_X1 U8748 ( .B1(n8084), .B2(n8087), .A(n15176), .ZN(n8082) );
  NAND2_X1 U8749 ( .A1(n15287), .A2(n8084), .ZN(n7702) );
  NOR2_X1 U8750 ( .A1(n13186), .A2(n15275), .ZN(n13196) );
  INV_X1 U8751 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n12183) );
  AND2_X1 U8752 ( .A1(n15235), .A2(n7693), .ZN(n7692) );
  INV_X1 U8753 ( .A(n15303), .ZN(n7693) );
  INV_X1 U8754 ( .A(n13210), .ZN(n13232) );
  NAND2_X1 U8755 ( .A1(n13232), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n13231) );
  NOR2_X1 U8756 ( .A1(n11305), .A2(n11304), .ZN(n11429) );
  OR2_X1 U8757 ( .A1(n11071), .A2(n11070), .ZN(n11305) );
  OR2_X1 U8758 ( .A1(n11969), .A2(n11968), .ZN(n12008) );
  OR2_X1 U8759 ( .A1(n11871), .A2(n12183), .ZN(n11969) );
  NAND2_X1 U8760 ( .A1(n11598), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n11871) );
  AND2_X1 U8761 ( .A1(n11429), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11598) );
  AND2_X1 U8762 ( .A1(n12056), .A2(n12054), .ZN(n7703) );
  NAND2_X1 U8763 ( .A1(n13302), .A2(n7666), .ZN(n13363) );
  NAND2_X1 U8764 ( .A1(n12990), .A2(n7667), .ZN(n7666) );
  INV_X1 U8765 ( .A(n13303), .ZN(n7667) );
  AND4_X1 U8766 ( .A1(n13010), .A2(n13009), .A3(n13008), .A4(n13007), .ZN(
        n15260) );
  AND4_X1 U8767 ( .A1(n13020), .A2(n13019), .A3(n13018), .A4(n13017), .ZN(
        n15636) );
  OR2_X1 U8768 ( .A1(n10529), .A2(n10349), .ZN(n10353) );
  NAND2_X1 U8769 ( .A1(n8317), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8314) );
  NOR2_X1 U8770 ( .A1(n15387), .A2(n15388), .ZN(n15386) );
  AOI21_X1 U8771 ( .B1(n15420), .B2(n10330), .A(n10329), .ZN(n10436) );
  AOI21_X1 U8772 ( .B1(n15451), .B2(n15450), .A(n15449), .ZN(n15448) );
  OR2_X1 U8773 ( .A1(n10210), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n10225) );
  OR2_X1 U8774 ( .A1(n10225), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n10232) );
  AOI21_X1 U8775 ( .B1(n11600), .B2(n10676), .A(n10675), .ZN(n10830) );
  XNOR2_X1 U8776 ( .A(n11483), .B(n12313), .ZN(n11485) );
  AOI21_X1 U8777 ( .B1(n12212), .B2(n12325), .A(n7584), .ZN(n12215) );
  AND2_X1 U8778 ( .A1(n12214), .A2(n12213), .ZN(n7584) );
  NAND2_X1 U8779 ( .A1(n15635), .A2(n8208), .ZN(n15607) );
  NAND2_X1 U8780 ( .A1(n7816), .A2(n7817), .ZN(n15612) );
  NAND2_X1 U8781 ( .A1(n15651), .A2(n7464), .ZN(n7816) );
  NAND2_X1 U8782 ( .A1(n15647), .A2(n7487), .ZN(n15629) );
  NAND2_X1 U8783 ( .A1(n15629), .A2(n15630), .ZN(n15628) );
  INV_X1 U8784 ( .A(n13231), .ZN(n13245) );
  NOR2_X1 U8785 ( .A1(n15676), .A2(n7785), .ZN(n7782) );
  INV_X1 U8786 ( .A(n8214), .ZN(n15665) );
  NOR2_X1 U8787 ( .A1(n15718), .A2(n15698), .ZN(n15701) );
  NAND2_X1 U8788 ( .A1(n15701), .A2(n15686), .ZN(n15685) );
  NAND2_X1 U8789 ( .A1(n8229), .A2(n8227), .ZN(n15680) );
  NAND2_X1 U8790 ( .A1(n13158), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13168) );
  OR2_X1 U8791 ( .A1(n13168), .A2(n13167), .ZN(n13186) );
  NOR2_X1 U8792 ( .A1(n15803), .A2(n15909), .ZN(n15792) );
  NAND2_X1 U8793 ( .A1(n15792), .A2(n15905), .ZN(n15774) );
  INV_X1 U8794 ( .A(n7870), .ZN(n7869) );
  AND2_X1 U8795 ( .A1(n7867), .A2(n8179), .ZN(n7866) );
  AOI21_X1 U8796 ( .B1(n8180), .B2(n8182), .A(n7504), .ZN(n8179) );
  NAND2_X1 U8797 ( .A1(n15568), .A2(n15567), .ZN(n15765) );
  NOR2_X1 U8798 ( .A1(n13122), .A2(n13121), .ZN(n13138) );
  NAND2_X1 U8799 ( .A1(n8216), .A2(n8215), .ZN(n15560) );
  AOI21_X1 U8800 ( .B1(n8217), .B2(n8219), .A(n7505), .ZN(n8215) );
  AND2_X1 U8801 ( .A1(n8235), .A2(n13324), .ZN(n8234) );
  OR2_X1 U8802 ( .A1(n8236), .A2(n7564), .ZN(n8235) );
  NAND2_X1 U8803 ( .A1(n11809), .A2(n8236), .ZN(n11870) );
  NOR2_X1 U8804 ( .A1(n11572), .A2(n8213), .ZN(n11816) );
  NOR2_X1 U8805 ( .A1(n11572), .A2(n16526), .ZN(n11815) );
  NOR2_X1 U8806 ( .A1(n11563), .A2(n8225), .ZN(n8224) );
  INV_X1 U8807 ( .A(n11567), .ZN(n8225) );
  NAND2_X1 U8808 ( .A1(n11059), .A2(n7447), .ZN(n8226) );
  NAND2_X1 U8809 ( .A1(n11211), .A2(n11216), .ZN(n11212) );
  INV_X1 U8810 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n10798) );
  NOR2_X1 U8811 ( .A1(n10799), .A2(n10798), .ZN(n10902) );
  NOR2_X1 U8812 ( .A1(n7865), .A2(n10869), .ZN(n7861) );
  INV_X1 U8813 ( .A(n10866), .ZN(n7865) );
  AND2_X1 U8814 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n10770) );
  INV_X1 U8815 ( .A(n15805), .ZN(n15787) );
  INV_X1 U8816 ( .A(n16389), .ZN(n15789) );
  INV_X1 U8817 ( .A(n7669), .ZN(n7668) );
  OAI22_X1 U8818 ( .A1(n7428), .A2(n7671), .B1(n13204), .B2(n7670), .ZN(n7669)
         );
  AND2_X1 U8819 ( .A1(n15253), .A2(n10871), .ZN(n11136) );
  INV_X1 U8820 ( .A(n10872), .ZN(n11122) );
  AND3_X1 U8821 ( .A1(n8211), .A2(n10470), .A3(n13308), .ZN(n11142) );
  NAND3_X1 U8822 ( .A1(n8315), .A2(n7449), .A3(n8316), .ZN(n13310) );
  NOR2_X1 U8823 ( .A1(n15582), .A2(n8200), .ZN(n8198) );
  INV_X1 U8824 ( .A(n15558), .ZN(n8200) );
  NAND2_X1 U8825 ( .A1(n8193), .A2(n15555), .ZN(n15688) );
  OR2_X1 U8826 ( .A1(n10407), .A2(n10409), .ZN(n16556) );
  XNOR2_X1 U8827 ( .A(n9310), .B(n9309), .ZN(n15104) );
  NAND2_X1 U8828 ( .A1(n10131), .A2(n8330), .ZN(n8329) );
  AND2_X1 U8829 ( .A1(n10220), .A2(n10217), .ZN(n8330) );
  INV_X1 U8830 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n10346) );
  XNOR2_X1 U8831 ( .A(n9338), .B(n9337), .ZN(n15112) );
  INV_X1 U8832 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10137) );
  XNOR2_X1 U8833 ( .A(n10216), .B(P1_IR_REG_21__SCAN_IN), .ZN(n12984) );
  NOR2_X1 U8834 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n8110) );
  XNOR2_X1 U8835 ( .A(n10358), .B(P1_IR_REG_19__SCAN_IN), .ZN(n13341) );
  NAND2_X1 U8836 ( .A1(n8257), .A2(n8487), .ZN(n8552) );
  OR2_X1 U8837 ( .A1(n8257), .A2(n7917), .ZN(n8905) );
  NAND2_X1 U8838 ( .A1(n8487), .A2(n8485), .ZN(n8903) );
  CLKBUF_X1 U8839 ( .A(n10123), .Z(n11009) );
  AND2_X1 U8840 ( .A1(n8870), .A2(n8869), .ZN(n13109) );
  NAND2_X1 U8841 ( .A1(n8278), .A2(n8476), .ZN(n8830) );
  NAND2_X1 U8842 ( .A1(n8280), .A2(n8279), .ZN(n8278) );
  INV_X1 U8843 ( .A(n8812), .ZN(n8280) );
  OR2_X1 U8844 ( .A1(n10384), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n10387) );
  OR2_X1 U8845 ( .A1(n10387), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n10648) );
  NAND2_X1 U8846 ( .A1(n7932), .A2(n8468), .ZN(n8770) );
  NAND2_X1 U8847 ( .A1(n8750), .A2(n8467), .ZN(n7932) );
  NAND2_X1 U8848 ( .A1(n8713), .A2(n8460), .ZN(n8731) );
  AOI21_X1 U8849 ( .B1(n8249), .B2(n8251), .A(n8248), .ZN(n8247) );
  INV_X1 U8850 ( .A(n8457), .ZN(n8248) );
  XNOR2_X1 U8851 ( .A(n8689), .B(n8688), .ZN(n11060) );
  NAND2_X1 U8852 ( .A1(n8674), .A2(n8452), .ZN(n8689) );
  OR2_X1 U8853 ( .A1(n10200), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n10189) );
  INV_X1 U8854 ( .A(SI_1_), .ZN(n7776) );
  INV_X1 U8855 ( .A(n8435), .ZN(n7777) );
  AND2_X1 U8856 ( .A1(n7891), .A2(n7889), .ZN(n16171) );
  NAND2_X1 U8857 ( .A1(n7890), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7889) );
  INV_X1 U8858 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7890) );
  OAI21_X1 U8859 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(n16217), .A(n16216), .ZN(
        n16225) );
  NAND2_X1 U8860 ( .A1(n16277), .A2(n16278), .ZN(n16290) );
  OAI22_X1 U8861 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n16302), .B1(n16301), 
        .B2(n16300), .ZN(n16307) );
  OR2_X1 U8862 ( .A1(n16339), .A2(n16338), .ZN(n16342) );
  XNOR2_X1 U8863 ( .A(n7705), .B(n13453), .ZN(n13454) );
  NAND2_X1 U8864 ( .A1(n13573), .A2(n13424), .ZN(n7705) );
  AND2_X1 U8865 ( .A1(n9795), .A2(n9794), .ZN(n13469) );
  INV_X1 U8866 ( .A(n13602), .ZN(n13807) );
  NOR2_X1 U8867 ( .A1(n13478), .A2(n13479), .ZN(n7722) );
  NAND2_X1 U8868 ( .A1(n13574), .A2(n13575), .ZN(n13573) );
  NAND2_X1 U8869 ( .A1(n7728), .A2(n7446), .ZN(n13406) );
  NAND2_X1 U8870 ( .A1(n13491), .A2(n8374), .ZN(n7728) );
  INV_X1 U8871 ( .A(n14001), .ZN(n13507) );
  AND2_X1 U8872 ( .A1(n9959), .A2(n9958), .ZN(n13779) );
  NAND2_X1 U8873 ( .A1(n8357), .A2(n8358), .ZN(n13510) );
  NAND2_X1 U8874 ( .A1(n13460), .A2(n8359), .ZN(n8357) );
  AND2_X1 U8875 ( .A1(n7720), .A2(n7721), .ZN(n12458) );
  INV_X1 U8876 ( .A(n13856), .ZN(n13879) );
  AND2_X1 U8877 ( .A1(n8378), .A2(n7481), .ZN(n13537) );
  NAND2_X1 U8878 ( .A1(n13491), .A2(n13490), .ZN(n8378) );
  INV_X1 U8879 ( .A(n13961), .ZN(n14055) );
  AND4_X1 U8880 ( .A1(n9801), .A2(n9800), .A3(n9799), .A4(n9798), .ZN(n13550)
         );
  NAND2_X1 U8881 ( .A1(n12616), .A2(n12615), .ZN(n12667) );
  NOR2_X1 U8882 ( .A1(n11193), .A2(n11192), .ZN(n11196) );
  INV_X1 U8883 ( .A(n7725), .ZN(n13480) );
  AND4_X1 U8884 ( .A1(n9851), .A2(n9850), .A3(n9849), .A4(n9848), .ZN(n13881)
         );
  NAND2_X1 U8885 ( .A1(n11040), .A2(n11039), .ZN(n13568) );
  INV_X1 U8886 ( .A(n13768), .ZN(n13733) );
  INV_X1 U8887 ( .A(n13599), .ZN(n13576) );
  AND2_X1 U8888 ( .A1(n10736), .A2(n11522), .ZN(n13596) );
  NAND2_X1 U8889 ( .A1(n13460), .A2(n8362), .ZN(n13584) );
  AND2_X1 U8890 ( .A1(n12743), .A2(n9585), .ZN(n13734) );
  INV_X1 U8891 ( .A(n13881), .ZN(n13904) );
  NAND4_X1 U8892 ( .A1(n9757), .A2(n9756), .A3(n9755), .A4(n9754), .ZN(n13953)
         );
  INV_X1 U8893 ( .A(n13971), .ZN(n12618) );
  NAND2_X1 U8894 ( .A1(n11090), .A2(n11089), .ZN(n11088) );
  XNOR2_X1 U8895 ( .A(n11721), .B(n11675), .ZN(n11664) );
  XNOR2_X1 U8896 ( .A(n11886), .B(n11893), .ZN(n11767) );
  INV_X1 U8897 ( .A(n7900), .ZN(n11887) );
  INV_X1 U8898 ( .A(n7899), .ZN(n11891) );
  INV_X1 U8899 ( .A(n7912), .ZN(n13642) );
  XNOR2_X1 U8900 ( .A(n7910), .B(n13668), .ZN(n13643) );
  NOR2_X1 U8901 ( .A1(n13643), .A2(n14037), .ZN(n13663) );
  INV_X1 U8902 ( .A(n13683), .ZN(n7638) );
  NOR2_X1 U8903 ( .A1(n10047), .A2(n10046), .ZN(n10048) );
  OR2_X1 U8904 ( .A1(n12733), .A2(n9644), .ZN(n9981) );
  NAND2_X1 U8905 ( .A1(n7627), .A2(n9595), .ZN(n9966) );
  NAND2_X1 U8906 ( .A1(n9927), .A2(n9926), .ZN(n13801) );
  NAND2_X1 U8907 ( .A1(n7986), .A2(n9915), .ZN(n13809) );
  NAND2_X1 U8908 ( .A1(n9908), .A2(n9907), .ZN(n14012) );
  NAND2_X1 U8909 ( .A1(n9884), .A2(n9883), .ZN(n14023) );
  OR2_X1 U8910 ( .A1(n10019), .A2(n7476), .ZN(n13865) );
  NAND2_X1 U8911 ( .A1(n7970), .A2(n12870), .ZN(n13863) );
  NAND2_X1 U8912 ( .A1(n13874), .A2(n13876), .ZN(n7970) );
  AND2_X1 U8913 ( .A1(n9830), .A2(n9829), .ZN(n13912) );
  NAND2_X1 U8914 ( .A1(n11522), .A2(n12920), .ZN(n13946) );
  NAND2_X1 U8915 ( .A1(n7962), .A2(n12829), .ZN(n12307) );
  NAND2_X1 U8916 ( .A1(n7607), .A2(n7444), .ZN(n7962) );
  OAI211_X1 U8917 ( .C1(SI_9_), .C2(n7430), .A(n9721), .B(n9720), .ZN(n12462)
         );
  INV_X1 U8918 ( .A(n13963), .ZN(n13942) );
  INV_X1 U8919 ( .A(n13977), .ZN(n13910) );
  NAND2_X1 U8920 ( .A1(n11521), .A2(n11520), .ZN(n13940) );
  INV_X1 U8921 ( .A(n13715), .ZN(n14067) );
  INV_X1 U8922 ( .A(n13720), .ZN(n14070) );
  AND3_X1 U8923 ( .A1(n13771), .A2(n13770), .A3(n13769), .ZN(n14079) );
  XNOR2_X1 U8924 ( .A(n13763), .B(n13764), .ZN(n14083) );
  XNOR2_X1 U8925 ( .A(n13777), .B(n13776), .ZN(n14089) );
  XNOR2_X1 U8926 ( .A(n13790), .B(n13791), .ZN(n14092) );
  AND2_X1 U8927 ( .A1(n9811), .A2(n9810), .ZN(n14123) );
  INV_X1 U8928 ( .A(n13469), .ZN(n14127) );
  NAND2_X1 U8929 ( .A1(n7607), .A2(n12825), .ZN(n12290) );
  OR2_X1 U8930 ( .A1(n10928), .A2(n10953), .ZN(n8017) );
  OR2_X1 U8931 ( .A1(n9644), .A2(n10144), .ZN(n8018) );
  AND2_X2 U8932 ( .A1(n10103), .A2(n10732), .ZN(n16590) );
  OR2_X1 U8933 ( .A1(n10237), .A2(P3_D_REG_1__SCAN_IN), .ZN(n10061) );
  NAND2_X1 U8934 ( .A1(n14140), .A2(n10237), .ZN(n10241) );
  NAND2_X1 U8935 ( .A1(n7620), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9553) );
  AOI21_X1 U8936 ( .B1(n9537), .B2(P1_DATAO_REG_24__SCAN_IN), .A(n9536), .ZN(
        n9934) );
  XNOR2_X1 U8937 ( .A(n9472), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12963) );
  INV_X1 U8938 ( .A(n12789), .ZN(n11442) );
  NAND2_X1 U8939 ( .A1(n8172), .A2(n7559), .ZN(n9896) );
  INV_X1 U8940 ( .A(SI_19_), .ZN(n14424) );
  INV_X1 U8941 ( .A(SI_18_), .ZN(n14425) );
  NAND2_X1 U8942 ( .A1(n8157), .A2(n8155), .ZN(n9856) );
  NAND2_X1 U8943 ( .A1(n8157), .A2(n7561), .ZN(n9854) );
  NAND2_X1 U8944 ( .A1(n9822), .A2(n9520), .ZN(n9839) );
  INV_X1 U8945 ( .A(SI_15_), .ZN(n14430) );
  INV_X1 U8946 ( .A(SI_14_), .ZN(n14435) );
  NAND2_X1 U8947 ( .A1(n7457), .A2(n8167), .ZN(n9775) );
  INV_X1 U8948 ( .A(SI_11_), .ZN(n14235) );
  INV_X1 U8949 ( .A(SI_10_), .ZN(n14440) );
  INV_X1 U8950 ( .A(SI_7_), .ZN(n10148) );
  INV_X1 U8951 ( .A(n8047), .ZN(n8046) );
  AND2_X1 U8952 ( .A1(n7629), .A2(n8705), .ZN(n8044) );
  NAND2_X1 U8953 ( .A1(n11460), .A2(n11461), .ZN(n11459) );
  NAND2_X1 U8954 ( .A1(n8940), .A2(n8939), .ZN(n15048) );
  NAND2_X1 U8955 ( .A1(n8666), .A2(n10722), .ZN(n10727) );
  NAND2_X1 U8956 ( .A1(n8897), .A2(n12537), .ZN(n12542) );
  NAND2_X1 U8957 ( .A1(n8021), .A2(n8995), .ZN(n14655) );
  NOR2_X1 U8958 ( .A1(n9441), .A2(n9405), .ZN(n8031) );
  INV_X1 U8959 ( .A(n10660), .ZN(n8032) );
  AOI21_X1 U8960 ( .B1(n8042), .B2(n8040), .A(n8039), .ZN(n8038) );
  INV_X1 U8961 ( .A(n8042), .ZN(n8041) );
  NAND2_X1 U8962 ( .A1(n11459), .A2(n8768), .ZN(n11693) );
  AOI21_X1 U8963 ( .B1(n10271), .B2(n10282), .A(n8117), .ZN(n8116) );
  NOR2_X1 U8964 ( .A1(n9357), .A2(n10172), .ZN(n8117) );
  NAND2_X1 U8965 ( .A1(n12542), .A2(n8901), .ZN(n14688) );
  NAND2_X1 U8966 ( .A1(n10727), .A2(n8670), .ZN(n11048) );
  AND2_X1 U8967 ( .A1(n8025), .A2(n8848), .ZN(n8024) );
  NAND2_X1 U8968 ( .A1(n9132), .A2(n14922), .ZN(n14691) );
  INV_X1 U8969 ( .A(n14700), .ZN(n14683) );
  NOR2_X1 U8970 ( .A1(n8431), .A2(n9450), .ZN(n9451) );
  NAND2_X1 U8971 ( .A1(n9342), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8575) );
  OR2_X1 U8972 ( .A1(n8969), .A2(n8579), .ZN(n8580) );
  OR2_X1 U8973 ( .A1(n8969), .A2(n10594), .ZN(n8596) );
  AND2_X1 U8974 ( .A1(n10312), .A2(P2_STATE_REG_SCAN_IN), .ZN(n16110) );
  INV_X1 U8975 ( .A(n14804), .ZN(n15000) );
  INV_X1 U8976 ( .A(n14810), .ZN(n15003) );
  AOI21_X1 U8977 ( .B1(n12696), .B2(n14981), .A(n12695), .ZN(n15009) );
  XNOR2_X1 U8978 ( .A(n7773), .B(n12716), .ZN(n12696) );
  NAND2_X1 U8979 ( .A1(n7743), .A2(n7440), .ZN(n14857) );
  NOR2_X1 U8980 ( .A1(n7490), .A2(n8058), .ZN(n14858) );
  NAND2_X1 U8981 ( .A1(n12686), .A2(n12685), .ZN(n14867) );
  NAND2_X1 U8982 ( .A1(n8131), .A2(n12709), .ZN(n14890) );
  NAND2_X1 U8983 ( .A1(n14899), .A2(n12708), .ZN(n8131) );
  NAND2_X1 U8984 ( .A1(n8964), .A2(n8963), .ZN(n15039) );
  OR2_X1 U8985 ( .A1(n12299), .A2(n9321), .ZN(n8964) );
  NAND2_X1 U8986 ( .A1(n12674), .A2(n12673), .ZN(n14979) );
  NAND2_X1 U8987 ( .A1(n8891), .A2(n8890), .ZN(n15068) );
  NAND2_X1 U8988 ( .A1(n12587), .A2(n12586), .ZN(n12588) );
  NAND2_X1 U8989 ( .A1(n12568), .A2(n12567), .ZN(n12570) );
  NAND2_X1 U8990 ( .A1(n12190), .A2(n12189), .ZN(n12262) );
  NAND2_X1 U8991 ( .A1(n8754), .A2(n8753), .ZN(n12151) );
  NAND2_X1 U8992 ( .A1(n12030), .A2(n11546), .ZN(n12070) );
  NAND2_X1 U8993 ( .A1(n8124), .A2(n11342), .ZN(n11919) );
  NAND2_X1 U8994 ( .A1(n8125), .A2(n7466), .ZN(n8124) );
  INV_X1 U8995 ( .A(n11341), .ZN(n8125) );
  NAND2_X2 U8996 ( .A1(n8657), .A2(n8656), .ZN(n11802) );
  NAND2_X1 U8997 ( .A1(n8063), .A2(n10818), .ZN(n10996) );
  INV_X1 U8998 ( .A(n8051), .ZN(n8050) );
  OAI22_X1 U8999 ( .A1(n9357), .A2(n10146), .B1(n8802), .B2(n16045), .ZN(n8051) );
  INV_X1 U9000 ( .A(n16515), .ZN(n16419) );
  INV_X1 U9001 ( .A(n7835), .ZN(n11323) );
  NAND2_X1 U9002 ( .A1(n10603), .A2(n10448), .ZN(n16622) );
  AND2_X1 U9003 ( .A1(n10270), .A2(P2_STATE_REG_SCAN_IN), .ZN(n16040) );
  OR2_X1 U9004 ( .A1(n15105), .A2(n8797), .ZN(n8540) );
  INV_X1 U9005 ( .A(n8508), .ZN(n8415) );
  XNOR2_X1 U9006 ( .A(n9106), .B(P2_IR_REG_26__SCAN_IN), .ZN(n15121) );
  NAND2_X1 U9007 ( .A1(n9110), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9106) );
  INV_X1 U9008 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12045) );
  NAND2_X1 U9009 ( .A1(n8529), .A2(n8515), .ZN(n8527) );
  INV_X1 U9010 ( .A(n9154), .ZN(n12727) );
  INV_X1 U9011 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10889) );
  INV_X1 U9012 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10643) );
  INV_X1 U9013 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10248) );
  OR2_X1 U9014 ( .A1(n8801), .A2(n8832), .ZN(n16126) );
  INV_X1 U9015 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10231) );
  INV_X1 U9016 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10229) );
  INV_X1 U9017 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10209) );
  INV_X1 U9018 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10173) );
  INV_X1 U9019 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10175) );
  INV_X1 U9020 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10160) );
  XNOR2_X1 U9021 ( .A(n10122), .B(n10121), .ZN(n10411) );
  NAND2_X1 U9022 ( .A1(n11109), .A2(n11108), .ZN(n11285) );
  NAND2_X1 U9023 ( .A1(n7698), .A2(n7697), .ZN(n11109) );
  NAND2_X1 U9024 ( .A1(n8093), .A2(n8098), .ZN(n15251) );
  NAND2_X1 U9025 ( .A1(n7688), .A2(n7451), .ZN(n8093) );
  NAND2_X1 U9026 ( .A1(n12516), .A2(n12515), .ZN(n12519) );
  NAND2_X1 U9027 ( .A1(n8115), .A2(n11613), .ZN(n11618) );
  NAND2_X1 U9028 ( .A1(n8091), .A2(n8094), .ZN(n15259) );
  AOI21_X1 U9029 ( .B1(n8098), .B2(n8100), .A(n15250), .ZN(n8094) );
  NOR2_X1 U9030 ( .A1(n8095), .A2(n7691), .ZN(n8092) );
  NAND2_X1 U9031 ( .A1(n8105), .A2(n11289), .ZN(n11302) );
  AND2_X1 U9032 ( .A1(n8114), .A2(n8113), .ZN(n15270) );
  AND2_X1 U9033 ( .A1(n12174), .A2(n12173), .ZN(n12181) );
  NAND2_X1 U9034 ( .A1(n10783), .A2(n7699), .ZN(n10890) );
  AOI21_X1 U9035 ( .B1(n15287), .B2(n15288), .A(n7439), .ZN(n15296) );
  INV_X1 U9036 ( .A(n7696), .ZN(n7686) );
  NAND2_X1 U9037 ( .A1(n15241), .A2(n15183), .ZN(n15310) );
  INV_X1 U9038 ( .A(n15876), .ZN(n15698) );
  NAND2_X1 U9039 ( .A1(n8083), .A2(n8088), .ZN(n15330) );
  NAND2_X1 U9040 ( .A1(n15287), .A2(n8089), .ZN(n8083) );
  NAND2_X1 U9041 ( .A1(n10527), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15360) );
  NAND2_X1 U9042 ( .A1(n7698), .A2(n10891), .ZN(n11104) );
  INV_X1 U9043 ( .A(n15367), .ZN(n15332) );
  NAND2_X1 U9044 ( .A1(n12405), .A2(n12404), .ZN(n15561) );
  NAND2_X1 U9045 ( .A1(n10425), .A2(n16395), .ZN(n15365) );
  OR2_X1 U9046 ( .A1(n13284), .A2(n16440), .ZN(n10484) );
  AOI21_X1 U9047 ( .B1(n11823), .B2(n10545), .A(n15474), .ZN(n15488) );
  XNOR2_X1 U9048 ( .A(n12214), .B(n12403), .ZN(n12212) );
  INV_X1 U9049 ( .A(n15526), .ZN(n15826) );
  NAND2_X1 U9050 ( .A1(n13292), .A2(n13291), .ZN(n15837) );
  NAND2_X1 U9051 ( .A1(n15600), .A2(n15599), .ZN(n15835) );
  AND2_X1 U9052 ( .A1(n13012), .A2(n13011), .ZN(n15621) );
  NAND2_X1 U9053 ( .A1(n15651), .A2(n15650), .ZN(n7818) );
  AND2_X1 U9054 ( .A1(n7878), .A2(n7877), .ZN(n15649) );
  NAND2_X1 U9055 ( .A1(n7783), .A2(n7784), .ZN(n15677) );
  NAND2_X1 U9056 ( .A1(n15866), .A2(n7879), .ZN(n15663) );
  NAND2_X1 U9057 ( .A1(n15996), .A2(n13204), .ZN(n15876) );
  NAND2_X1 U9058 ( .A1(n15716), .A2(n8232), .ZN(n15695) );
  AND2_X1 U9059 ( .A1(n15716), .A2(n15574), .ZN(n15697) );
  INV_X1 U9060 ( .A(n8228), .ZN(n8232) );
  INV_X1 U9061 ( .A(n15724), .ZN(n15552) );
  NAND2_X1 U9062 ( .A1(n8190), .A2(n15548), .ZN(n15742) );
  NAND2_X1 U9063 ( .A1(n13179), .A2(n13178), .ZN(n15889) );
  NAND2_X1 U9064 ( .A1(n15767), .A2(n15569), .ZN(n15751) );
  NAND2_X1 U9065 ( .A1(n15815), .A2(n15543), .ZN(n15784) );
  NAND2_X1 U9066 ( .A1(n12317), .A2(n12316), .ZN(n12319) );
  NAND2_X1 U9067 ( .A1(n12311), .A2(n12310), .ZN(n12409) );
  NAND2_X1 U9068 ( .A1(n11962), .A2(n11961), .ZN(n13090) );
  NAND2_X1 U9069 ( .A1(n11861), .A2(n11860), .ZN(n11866) );
  AND2_X1 U9070 ( .A1(n11809), .A2(n11593), .ZN(n11594) );
  NAND2_X1 U9071 ( .A1(n11583), .A2(n11582), .ZN(n11808) );
  NAND2_X1 U9072 ( .A1(n11562), .A2(n11561), .ZN(n11564) );
  NAND2_X1 U9073 ( .A1(n11059), .A2(n11058), .ZN(n11568) );
  NAND2_X1 U9074 ( .A1(n10867), .A2(n10866), .ZN(n11370) );
  INV_X1 U9075 ( .A(n15780), .ZN(n16601) );
  NAND2_X1 U9076 ( .A1(n15812), .A2(n11128), .ZN(n16595) );
  NAND2_X1 U9077 ( .A1(n10494), .A2(n13289), .ZN(n7860) );
  INV_X1 U9078 ( .A(n7859), .ZN(n7858) );
  AND2_X1 U9079 ( .A1(n15812), .A2(n16458), .ZN(n15711) );
  NAND2_X1 U9080 ( .A1(n15812), .A2(n11136), .ZN(n16597) );
  INV_X1 U9081 ( .A(n16595), .ZN(n16525) );
  OAI211_X1 U9082 ( .C1(n15838), .C2(n16435), .A(n7804), .B(n7602), .ZN(n15948) );
  NOR2_X1 U9083 ( .A1(n15836), .A2(n7805), .ZN(n7804) );
  INV_X1 U9084 ( .A(n15835), .ZN(n7602) );
  AND2_X1 U9085 ( .A1(n15837), .A2(n16490), .ZN(n7805) );
  AND2_X1 U9086 ( .A1(n10133), .A2(n10219), .ZN(n10391) );
  NAND2_X1 U9087 ( .A1(n9319), .A2(n9320), .ZN(n15975) );
  INV_X1 U9088 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10342) );
  INV_X1 U9089 ( .A(n10391), .ZN(n15985) );
  NAND2_X1 U9090 ( .A1(n7701), .A2(n7700), .ZN(n10136) );
  NAND2_X1 U9091 ( .A1(n10130), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7700) );
  OAI21_X1 U9092 ( .B1(n10134), .B2(n10344), .A(P1_IR_REG_25__SCAN_IN), .ZN(
        n7701) );
  NAND2_X1 U9093 ( .A1(n8983), .A2(n8982), .ZN(n8997) );
  XNOR2_X1 U9094 ( .A(n7939), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15996) );
  NAND2_X1 U9095 ( .A1(n13203), .A2(n10165), .ZN(n7939) );
  INV_X1 U9096 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n13177) );
  INV_X1 U9097 ( .A(n13341), .ZN(n15519) );
  INV_X1 U9098 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11473) );
  INV_X1 U9099 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11244) );
  NAND2_X1 U9100 ( .A1(n7652), .A2(n10115), .ZN(n11242) );
  INV_X1 U9101 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10650) );
  INV_X1 U9102 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10601) );
  INV_X1 U9103 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10252) );
  INV_X1 U9104 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10235) );
  INV_X1 U9105 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10227) );
  INV_X1 U9106 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10205) );
  INV_X1 U9107 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10192) );
  NAND2_X1 U9108 ( .A1(n8673), .A2(n8674), .ZN(n10892) );
  INV_X1 U9109 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10195) );
  INV_X1 U9110 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10186) );
  MUX2_X1 U9111 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10169), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n10171) );
  INV_X1 U9112 ( .A(P2_RD_REG_SCAN_IN), .ZN(n16385) );
  NAND2_X1 U9113 ( .A1(n16221), .A2(n7894), .ZN(n16354) );
  INV_X1 U9114 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7895) );
  NOR2_X1 U9115 ( .A1(n16272), .A2(n16273), .ZN(n16274) );
  XNOR2_X1 U9116 ( .A(n16290), .B(n7888), .ZN(n16284) );
  INV_X1 U9117 ( .A(n16291), .ZN(n7888) );
  NAND2_X1 U9118 ( .A1(n12157), .A2(n12156), .ZN(n12159) );
  INV_X1 U9119 ( .A(n7909), .ZN(n12487) );
  INV_X1 U9120 ( .A(n7737), .ZN(n12491) );
  NAND2_X1 U9121 ( .A1(n9128), .A2(n14707), .ZN(n9153) );
  NAND2_X1 U9122 ( .A1(n8023), .A2(n12132), .ZN(n12138) );
  AOI21_X1 U9123 ( .B1(n14193), .B2(n7474), .A(n7631), .ZN(n14198) );
  NAND2_X1 U9124 ( .A1(n14195), .A2(n7632), .ZN(n7631) );
  AOI211_X1 U9125 ( .C1(n16508), .C2(n15010), .A(n14831), .B(n14830), .ZN(
        n14832) );
  INV_X1 U9126 ( .A(n7660), .ZN(n13370) );
  OR2_X1 U9127 ( .A1(n16469), .A2(n13006), .ZN(n7933) );
  NAND2_X1 U9128 ( .A1(n7882), .A2(n16469), .ZN(n7934) );
  NAND2_X1 U9129 ( .A1(n16564), .A2(n16570), .ZN(n8197) );
  INV_X1 U9130 ( .A(n8196), .ZN(n8195) );
  OAI21_X1 U9131 ( .B1(n15833), .B2(n16567), .A(n8202), .ZN(n8196) );
  NAND2_X1 U9132 ( .A1(n7803), .A2(n7802), .ZN(P1_U3524) );
  NAND2_X1 U9133 ( .A1(n16567), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7802) );
  NAND2_X1 U9134 ( .A1(n15948), .A2(n16570), .ZN(n7803) );
  NAND2_X1 U9135 ( .A1(n15949), .A2(n16570), .ZN(n8240) );
  INV_X1 U9136 ( .A(n16245), .ZN(n16241) );
  XNOR2_X1 U9137 ( .A(n7885), .B(n7630), .ZN(SUB_1596_U4) );
  XNOR2_X1 U9138 ( .A(n16352), .B(n16351), .ZN(n7630) );
  NAND2_X1 U9139 ( .A1(n16348), .A2(n7886), .ZN(n7885) );
  AND4_X1 U9140 ( .A1(n8430), .A2(n8507), .A3(n8516), .A4(n8528), .ZN(n7438)
         );
  INV_X1 U9141 ( .A(n14822), .ZN(n8078) );
  INV_X2 U9142 ( .A(n10797), .ZN(n13277) );
  NAND2_X1 U9143 ( .A1(n13439), .A2(n9580), .ZN(n9649) );
  INV_X2 U9144 ( .A(n9649), .ZN(n10038) );
  INV_X2 U9145 ( .A(n9649), .ZN(n9984) );
  AND2_X1 U9146 ( .A1(n15162), .A2(n15161), .ZN(n7439) );
  INV_X1 U9147 ( .A(n15281), .ZN(n7691) );
  AND2_X1 U9148 ( .A1(n7517), .A2(n7747), .ZN(n7440) );
  INV_X1 U9149 ( .A(n15383), .ZN(n7856) );
  NAND2_X1 U9150 ( .A1(n9579), .A2(n9580), .ZN(n9662) );
  AND2_X1 U9151 ( .A1(n7709), .A2(n13526), .ZN(n7441) );
  OR2_X1 U9152 ( .A1(n8483), .A2(SI_17_), .ZN(n7442) );
  AND2_X1 U9153 ( .A1(n7966), .A2(n12825), .ZN(n7444) );
  INV_X1 U9154 ( .A(n12706), .ZN(n7770) );
  AND2_X1 U9155 ( .A1(n15687), .A2(n8227), .ZN(n7445) );
  AND2_X1 U9156 ( .A1(n8377), .A2(n13393), .ZN(n7446) );
  AND2_X1 U9157 ( .A1(n7484), .A2(n11058), .ZN(n7447) );
  AND2_X1 U9158 ( .A1(n8343), .A2(n12666), .ZN(n7448) );
  AND2_X1 U9159 ( .A1(n10354), .A2(n10352), .ZN(n7449) );
  AND2_X1 U9160 ( .A1(n12675), .A2(n7761), .ZN(n7450) );
  INV_X1 U9161 ( .A(n11173), .ZN(n16452) );
  INV_X1 U9162 ( .A(n9245), .ZN(n8420) );
  INV_X1 U9163 ( .A(n11754), .ZN(n12163) );
  NOR2_X1 U9164 ( .A1(n7690), .A2(n8100), .ZN(n7451) );
  AOI21_X1 U9165 ( .B1(n9288), .B2(n7548), .A(n7855), .ZN(n9290) );
  AND2_X1 U9166 ( .A1(n13002), .A2(n13001), .ZN(n15830) );
  AND2_X1 U9167 ( .A1(n7521), .A2(n8420), .ZN(n7452) );
  AND2_X1 U9168 ( .A1(n8118), .A2(n12592), .ZN(n7453) );
  INV_X1 U9169 ( .A(n14821), .ZN(n8076) );
  NAND2_X1 U9170 ( .A1(n8360), .A2(n8363), .ZN(n8359) );
  INV_X1 U9171 ( .A(n8359), .ZN(n8353) );
  NAND2_X1 U9172 ( .A1(n8324), .A2(n8325), .ZN(n7454) );
  AND4_X1 U9173 ( .A1(n10127), .A2(n10126), .A3(n10125), .A4(n10124), .ZN(
        n7455) );
  NAND3_X1 U9174 ( .A1(n8516), .A2(n8906), .A3(n8515), .ZN(n7456) );
  INV_X1 U9175 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n10116) );
  INV_X1 U9176 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n9556) );
  NAND2_X1 U9177 ( .A1(n12806), .A2(n9647), .ZN(n9995) );
  INV_X1 U9178 ( .A(n9995), .ZN(n7578) );
  AND2_X1 U9179 ( .A1(n8168), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7457) );
  INV_X1 U9180 ( .A(n13180), .ZN(n7684) );
  AND2_X1 U9181 ( .A1(n8416), .A2(n8542), .ZN(n7458) );
  NAND2_X1 U9182 ( .A1(n13295), .A2(n8323), .ZN(n7459) );
  INV_X1 U9183 ( .A(n9159), .ZN(n9168) );
  AND2_X1 U9184 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n9514), .ZN(n7460) );
  NAND2_X1 U9185 ( .A1(n7725), .A2(n7722), .ZN(n7727) );
  NAND2_X1 U9186 ( .A1(n11928), .A2(n16516), .ZN(n12035) );
  INV_X1 U9187 ( .A(n12035), .ZN(n7948) );
  NAND2_X1 U9188 ( .A1(n10348), .A2(n15979), .ZN(n10797) );
  NOR2_X1 U9189 ( .A1(n12289), .A2(n12828), .ZN(n7461) );
  NAND2_X1 U9190 ( .A1(n8161), .A2(n10389), .ZN(n8167) );
  OAI211_X1 U9191 ( .C1(n9645), .C2(SI_4_), .A(n8018), .B(n8017), .ZN(n8016)
         );
  AND2_X1 U9192 ( .A1(n9002), .A2(n9001), .ZN(n14889) );
  INV_X1 U9193 ( .A(n14889), .ZN(n15030) );
  OR4_X1 U9194 ( .A1(n13340), .A2(n13000), .A3(n13347), .A4(n13358), .ZN(n7463) );
  NAND2_X1 U9195 ( .A1(n15241), .A2(n8111), .ZN(n8114) );
  NAND2_X1 U9196 ( .A1(n8345), .A2(n8347), .ZN(n10053) );
  AND2_X1 U9197 ( .A1(n7822), .A2(n15650), .ZN(n7464) );
  XOR2_X1 U9198 ( .A(n14012), .B(n13428), .Z(n7465) );
  AOI21_X1 U9199 ( .B1(n8331), .B2(n13526), .A(n7711), .ZN(n7710) );
  OR2_X1 U9200 ( .A1(n11802), .A2(n14731), .ZN(n7466) );
  INV_X1 U9201 ( .A(n15979), .ZN(n10350) );
  OR2_X1 U9202 ( .A1(n9178), .A2(n9177), .ZN(n7467) );
  INV_X1 U9203 ( .A(n13508), .ZN(n8356) );
  NOR2_X2 U9204 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8570) );
  NAND3_X1 U9205 ( .A1(n8345), .A2(n8347), .A3(n7987), .ZN(n7468) );
  NOR2_X1 U9206 ( .A1(n13660), .A2(n7642), .ZN(n7469) );
  AND2_X1 U9207 ( .A1(n12898), .A2(n12899), .ZN(n7470) );
  AND2_X1 U9208 ( .A1(n7694), .A2(n7695), .ZN(n7471) );
  AND2_X1 U9209 ( .A1(n8290), .A2(n7658), .ZN(n7472) );
  XNOR2_X1 U9210 ( .A(n10215), .B(n10214), .ZN(n12983) );
  NOR2_X1 U9211 ( .A1(n9624), .A2(n8367), .ZN(n9641) );
  OR2_X1 U9212 ( .A1(n8620), .A2(n10280), .ZN(n7473) );
  AND3_X1 U9213 ( .A1(n14199), .A2(n14192), .A3(n14707), .ZN(n7474) );
  NAND2_X1 U9214 ( .A1(n15380), .A2(n13053), .ZN(n7475) );
  AND2_X1 U9215 ( .A1(n13884), .A2(n13868), .ZN(n7476) );
  OR3_X1 U9216 ( .A1(n9388), .A2(n9387), .A3(n9386), .ZN(n7477) );
  INV_X1 U9217 ( .A(n10123), .ZN(n7652) );
  NOR2_X1 U9218 ( .A1(n14012), .A2(n13833), .ZN(n7478) );
  NAND2_X1 U9219 ( .A1(n13252), .A2(n13251), .ZN(n15853) );
  NAND2_X1 U9220 ( .A1(n9074), .A2(n9073), .ZN(n14843) );
  AND3_X1 U9221 ( .A1(n12955), .A2(n13694), .A3(n12957), .ZN(n7479) );
  NAND2_X1 U9222 ( .A1(n13413), .A2(n13526), .ZN(n13472) );
  AND2_X1 U9223 ( .A1(n8052), .A2(n12594), .ZN(n7480) );
  OR2_X1 U9224 ( .A1(n13390), .A2(n13879), .ZN(n7481) );
  AND2_X1 U9225 ( .A1(n15281), .A2(n7692), .ZN(n7482) );
  AND2_X1 U9226 ( .A1(n15847), .A2(n15653), .ZN(n7483) );
  OR2_X1 U9227 ( .A1(n13065), .A2(n11566), .ZN(n7484) );
  NAND2_X1 U9228 ( .A1(n11418), .A2(n11417), .ZN(n13078) );
  NAND2_X1 U9229 ( .A1(n13413), .A2(n13824), .ZN(n8331) );
  INV_X1 U9230 ( .A(n8331), .ZN(n7709) );
  AND2_X1 U9231 ( .A1(n15271), .A2(n8113), .ZN(n7485) );
  INV_X1 U9232 ( .A(n7427), .ZN(n14852) );
  NOR3_X1 U9233 ( .A1(n14918), .A2(n7949), .A3(n15022), .ZN(n7604) );
  AND2_X1 U9234 ( .A1(n12095), .A2(n14727), .ZN(n7486) );
  NAND2_X1 U9235 ( .A1(n13239), .A2(n13238), .ZN(n15859) );
  INV_X1 U9236 ( .A(n9253), .ZN(n8414) );
  NAND2_X1 U9237 ( .A1(n8346), .A2(n8347), .ZN(n10051) );
  OR2_X1 U9238 ( .A1(n15655), .A2(n15579), .ZN(n7487) );
  OR2_X1 U9239 ( .A1(n11893), .A2(n11886), .ZN(n7488) );
  AND2_X1 U9240 ( .A1(n7640), .A2(n7639), .ZN(n7489) );
  AND2_X1 U9241 ( .A1(n9051), .A2(n9050), .ZN(n14856) );
  INV_X1 U9242 ( .A(n14856), .ZN(n15022) );
  INV_X1 U9243 ( .A(n8276), .ZN(n8275) );
  NOR2_X1 U9244 ( .A1(n8829), .A2(n8277), .ZN(n8276) );
  NAND2_X1 U9245 ( .A1(n8835), .A2(n8834), .ZN(n12566) );
  AND2_X1 U9246 ( .A1(n12686), .A2(n8056), .ZN(n7490) );
  INV_X1 U9247 ( .A(n7880), .ZN(n7879) );
  INV_X2 U9248 ( .A(n12736), .ZN(n10039) );
  INV_X1 U9249 ( .A(n8363), .ZN(n8362) );
  NAND2_X1 U9250 ( .A1(n13953), .A2(n14060), .ZN(n7491) );
  AND2_X1 U9251 ( .A1(n9029), .A2(n9028), .ZN(n14877) );
  INV_X1 U9252 ( .A(n14877), .ZN(n7953) );
  AND2_X1 U9253 ( .A1(n8131), .A2(n8129), .ZN(n7492) );
  OR2_X1 U9254 ( .A1(n12486), .A2(n12485), .ZN(n7493) );
  AND2_X1 U9255 ( .A1(n8322), .A2(n7459), .ZN(n7494) );
  AND2_X1 U9256 ( .A1(n14889), .A2(n14870), .ZN(n7495) );
  AND2_X1 U9257 ( .A1(n10033), .A2(n10032), .ZN(n7496) );
  AND2_X1 U9258 ( .A1(n12517), .A2(n12515), .ZN(n7497) );
  AND2_X1 U9259 ( .A1(n14843), .A2(n14861), .ZN(n7498) );
  NAND2_X1 U9260 ( .A1(n14031), .A2(n13868), .ZN(n12870) );
  INV_X1 U9261 ( .A(n12870), .ZN(n7973) );
  AND2_X1 U9262 ( .A1(n13811), .A2(n13794), .ZN(n7499) );
  INV_X1 U9263 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8542) );
  AND2_X1 U9264 ( .A1(n16499), .A2(n11350), .ZN(n7500) );
  AND2_X1 U9265 ( .A1(n8327), .A2(n10346), .ZN(n7501) );
  AND2_X1 U9266 ( .A1(n14995), .A2(n14718), .ZN(n7502) );
  NOR2_X1 U9267 ( .A1(n14877), .A2(n14860), .ZN(n7503) );
  OR2_X1 U9268 ( .A1(n7778), .A2(n10164), .ZN(n7755) );
  NOR2_X1 U9269 ( .A1(n15909), .A2(n15768), .ZN(n7504) );
  NOR2_X1 U9270 ( .A1(n13102), .A2(n15358), .ZN(n7505) );
  AND2_X1 U9271 ( .A1(n8412), .A2(n9253), .ZN(n7506) );
  AND2_X1 U9272 ( .A1(n12618), .A2(n12617), .ZN(n7507) );
  OR2_X1 U9273 ( .A1(n7684), .A2(n7683), .ZN(n7508) );
  INV_X1 U9274 ( .A(n7785), .ZN(n7784) );
  NOR2_X1 U9275 ( .A1(n15686), .A2(n15703), .ZN(n7785) );
  NAND2_X1 U9276 ( .A1(n10470), .A2(n8211), .ZN(n13025) );
  INV_X1 U9277 ( .A(n8183), .ZN(n7877) );
  NOR2_X1 U9278 ( .A1(n15859), .A2(n15577), .ZN(n8183) );
  INV_X1 U9279 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7671) );
  NAND2_X1 U9280 ( .A1(n7778), .A2(n7750), .ZN(n7509) );
  AND2_X1 U9281 ( .A1(n8392), .A2(n7623), .ZN(n7510) );
  NAND2_X1 U9282 ( .A1(n8172), .A2(n9526), .ZN(n7511) );
  INV_X1 U9283 ( .A(n8209), .ZN(n8208) );
  NAND2_X1 U9284 ( .A1(n15621), .A2(n8210), .ZN(n8209) );
  INV_X1 U9285 ( .A(n7999), .ZN(n7998) );
  AND2_X1 U9286 ( .A1(n13808), .A2(n8000), .ZN(n7999) );
  AND2_X1 U9287 ( .A1(n8479), .A2(n14430), .ZN(n7512) );
  INV_X1 U9288 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n9657) );
  INV_X1 U9289 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8514) );
  NAND2_X1 U9290 ( .A1(n9268), .A2(n9269), .ZN(n7513) );
  NOR2_X1 U9291 ( .A1(n12954), .A2(n12953), .ZN(n7514) );
  AND2_X1 U9292 ( .A1(n8478), .A2(n14435), .ZN(n7515) );
  AND2_X1 U9293 ( .A1(n8470), .A2(n14235), .ZN(n7516) );
  AND2_X1 U9294 ( .A1(n14859), .A2(n12687), .ZN(n7517) );
  AND2_X1 U9295 ( .A1(n8787), .A2(n8786), .ZN(n7518) );
  INV_X1 U9296 ( .A(n15598), .ZN(n7811) );
  AND2_X1 U9297 ( .A1(n12690), .A2(n9417), .ZN(n14822) );
  OR2_X1 U9298 ( .A1(n7430), .A2(SI_3_), .ZN(n7519) );
  AND2_X1 U9299 ( .A1(n7771), .A2(n12680), .ZN(n7520) );
  AND2_X1 U9300 ( .A1(n9244), .A2(n9243), .ZN(n7521) );
  AND2_X1 U9301 ( .A1(n9157), .A2(n9405), .ZN(n7522) );
  INV_X1 U9302 ( .A(n7820), .ZN(n7814) );
  NAND2_X1 U9303 ( .A1(n15840), .A2(n15636), .ZN(n7820) );
  NAND2_X1 U9304 ( .A1(n7524), .A2(n7822), .ZN(n7817) );
  NAND2_X1 U9305 ( .A1(n8324), .A2(n13276), .ZN(n7523) );
  INV_X1 U9306 ( .A(n13083), .ZN(n7659) );
  INV_X1 U9307 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n10130) );
  INV_X1 U9308 ( .A(n8395), .ZN(n8394) );
  NAND2_X1 U9309 ( .A1(n9218), .A2(n9220), .ZN(n8395) );
  OR2_X1 U9310 ( .A1(n7819), .A2(n7483), .ZN(n7524) );
  INV_X1 U9311 ( .A(n13181), .ZN(n7681) );
  INV_X1 U9312 ( .A(n13240), .ZN(n7677) );
  INV_X1 U9313 ( .A(n13308), .ZN(n8315) );
  INV_X1 U9314 ( .A(n15547), .ZN(n15757) );
  NAND2_X1 U9315 ( .A1(n11587), .A2(n11586), .ZN(n13082) );
  NOR2_X1 U9316 ( .A1(n13405), .A2(n7465), .ZN(n7525) );
  NAND4_X1 U9317 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n10483), .ZN(
        n15383) );
  AND2_X1 U9318 ( .A1(n13402), .A2(n10021), .ZN(n13835) );
  INV_X1 U9319 ( .A(n13835), .ZN(n7581) );
  OR2_X1 U9320 ( .A1(n8350), .A2(n8352), .ZN(n7526) );
  AND2_X1 U9321 ( .A1(n12650), .A2(n12648), .ZN(n7527) );
  AND2_X1 U9322 ( .A1(n10029), .A2(n12768), .ZN(n13777) );
  AND2_X1 U9323 ( .A1(n10868), .A2(n7475), .ZN(n7528) );
  AND2_X1 U9324 ( .A1(n11620), .A2(n11613), .ZN(n7529) );
  NOR2_X1 U9325 ( .A1(n8123), .A2(n11918), .ZN(n8122) );
  NOR2_X1 U9326 ( .A1(n7790), .A2(n7929), .ZN(n7789) );
  NAND2_X1 U9327 ( .A1(n11105), .A2(n11103), .ZN(n7530) );
  AND2_X1 U9328 ( .A1(n7713), .A2(n8342), .ZN(n7531) );
  AND2_X1 U9329 ( .A1(n10009), .A2(n8006), .ZN(n7532) );
  AND2_X1 U9330 ( .A1(n7740), .A2(n8449), .ZN(n7533) );
  AND2_X1 U9331 ( .A1(n8147), .A2(n9540), .ZN(n7534) );
  NAND2_X1 U9332 ( .A1(n13088), .A2(n8296), .ZN(n7535) );
  OR2_X1 U9333 ( .A1(n7506), .A2(n7838), .ZN(n7536) );
  AND2_X1 U9334 ( .A1(n8310), .A2(n7676), .ZN(n7537) );
  AND2_X1 U9335 ( .A1(n8306), .A2(n7682), .ZN(n7538) );
  NAND2_X1 U9336 ( .A1(n13133), .A2(n8305), .ZN(n7539) );
  NAND2_X1 U9337 ( .A1(n13100), .A2(n8299), .ZN(n7540) );
  AND2_X1 U9338 ( .A1(n9181), .A2(n9180), .ZN(n7541) );
  INV_X1 U9339 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n10217) );
  NAND2_X1 U9340 ( .A1(n15341), .A2(n8101), .ZN(n8100) );
  NAND2_X1 U9341 ( .A1(n13107), .A2(n8302), .ZN(n7542) );
  INV_X1 U9342 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n14143) );
  INV_X1 U9343 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10146) );
  INV_X1 U9344 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10164) );
  INV_X1 U9345 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10172) );
  INV_X1 U9346 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8509) );
  INV_X1 U9347 ( .A(n8135), .ZN(n8134) );
  NAND2_X1 U9348 ( .A1(n12715), .A2(n8136), .ZN(n8135) );
  OR2_X1 U9349 ( .A1(n13994), .A2(n13993), .ZN(P3_U3486) );
  OR2_X1 U9350 ( .A1(n14078), .A2(n14077), .ZN(P3_U3454) );
  OR2_X1 U9351 ( .A1(n13762), .A2(n13761), .ZN(P3_U3206) );
  INV_X1 U9352 ( .A(n14992), .ZN(n14954) );
  AND2_X2 U9353 ( .A1(n11787), .A2(n14922), .ZN(n14992) );
  INV_X1 U9354 ( .A(n11385), .ZN(n7908) );
  INV_X1 U9355 ( .A(n13817), .ZN(n7982) );
  INV_X1 U9356 ( .A(n15726), .ZN(n7873) );
  INV_X1 U9357 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8109) );
  INV_X1 U9358 ( .A(n14967), .ZN(n7583) );
  NAND2_X1 U9359 ( .A1(n8985), .A2(n8984), .ZN(n15035) );
  INV_X1 U9360 ( .A(n15035), .ZN(n7952) );
  NAND2_X1 U9361 ( .A1(n12193), .A2(n12194), .ZN(n12266) );
  INV_X1 U9362 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10389) );
  INV_X1 U9363 ( .A(n13284), .ZN(n8317) );
  INV_X1 U9364 ( .A(n8811), .ZN(n8279) );
  INV_X1 U9365 ( .A(n12828), .ZN(n7966) );
  NAND2_X1 U9366 ( .A1(n12302), .A2(n10007), .ZN(n12475) );
  NAND2_X1 U9367 ( .A1(n12879), .A2(n12880), .ZN(n13852) );
  INV_X1 U9368 ( .A(n13852), .ZN(n7579) );
  AND2_X1 U9369 ( .A1(n15614), .A2(n15787), .ZN(n7546) );
  AND2_X1 U9370 ( .A1(n12593), .A2(n12592), .ZN(n7547) );
  AND2_X1 U9371 ( .A1(n9286), .A2(n9285), .ZN(n7548) );
  AND2_X1 U9372 ( .A1(n15621), .A2(n15636), .ZN(n7549) );
  OR2_X1 U9373 ( .A1(n7851), .A2(n7847), .ZN(n7550) );
  NAND2_X1 U9374 ( .A1(n7848), .A2(n7846), .ZN(n7551) );
  AND2_X1 U9375 ( .A1(n9252), .A2(n9251), .ZN(n7552) );
  INV_X1 U9376 ( .A(n8902), .ZN(n8486) );
  INV_X1 U9377 ( .A(n7597), .ZN(n15802) );
  NOR2_X1 U9378 ( .A1(n12410), .A2(n15561), .ZN(n7597) );
  AND2_X1 U9379 ( .A1(n8959), .A2(SI_21_), .ZN(n7553) );
  NAND2_X1 U9380 ( .A1(n9950), .A2(n9949), .ZN(n8177) );
  INV_X1 U9381 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10492) );
  OR2_X1 U9382 ( .A1(n12503), .A2(n12500), .ZN(n7554) );
  AND2_X1 U9383 ( .A1(n12173), .A2(n12180), .ZN(n7555) );
  AND2_X1 U9384 ( .A1(n12055), .A2(n12054), .ZN(n7556) );
  AND2_X1 U9385 ( .A1(n12649), .A2(n12648), .ZN(n7557) );
  AND2_X1 U9386 ( .A1(n12072), .A2(n12071), .ZN(n7558) );
  INV_X1 U9387 ( .A(n7923), .ZN(n7922) );
  NOR2_X1 U9388 ( .A1(n8284), .A2(n7924), .ZN(n7923) );
  INV_X1 U9389 ( .A(n7821), .ZN(n7819) );
  NAND2_X1 U9390 ( .A1(n15853), .A2(n15579), .ZN(n7821) );
  INV_X1 U9391 ( .A(n7442), .ZN(n7799) );
  INV_X1 U9392 ( .A(n12594), .ZN(n8118) );
  INV_X1 U9393 ( .A(n12132), .ZN(n8027) );
  AND2_X1 U9394 ( .A1(n9893), .A2(n9526), .ZN(n7559) );
  NAND2_X1 U9395 ( .A1(n13112), .A2(n13111), .ZN(n15919) );
  INV_X1 U9396 ( .A(n15919), .ZN(n7596) );
  INV_X1 U9397 ( .A(n12537), .ZN(n8040) );
  NAND2_X2 U9398 ( .A1(n12963), .A2(n12789), .ZN(n12901) );
  AND2_X1 U9399 ( .A1(n12078), .A2(n7954), .ZN(n7560) );
  OR2_X1 U9400 ( .A1(n11244), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7561) );
  INV_X1 U9401 ( .A(n11572), .ZN(n7599) );
  NAND2_X1 U9402 ( .A1(n11748), .A2(n12816), .ZN(n12106) );
  NAND2_X1 U9403 ( .A1(n7864), .A2(n10868), .ZN(n11064) );
  NOR2_X1 U9404 ( .A1(n8519), .A2(n9405), .ZN(n9130) );
  INV_X1 U9405 ( .A(n8960), .ZN(n8256) );
  AND2_X1 U9406 ( .A1(n15168), .A2(n15167), .ZN(n7562) );
  OR2_X1 U9407 ( .A1(n11572), .A2(n8212), .ZN(n7563) );
  NOR2_X1 U9408 ( .A1(n13082), .A2(n11868), .ZN(n7564) );
  NAND2_X1 U9409 ( .A1(n8003), .A2(n10001), .ZN(n12241) );
  AND2_X1 U9410 ( .A1(n7727), .A2(n8332), .ZN(n7565) );
  AND2_X1 U9411 ( .A1(n8226), .A2(n8224), .ZN(n7566) );
  AND2_X1 U9412 ( .A1(n8066), .A2(n8067), .ZN(n7567) );
  NAND2_X1 U9413 ( .A1(n10792), .A2(n10793), .ZN(n7568) );
  INV_X1 U9414 ( .A(n8156), .ZN(n8155) );
  NAND2_X1 U9415 ( .A1(n8160), .A2(n7561), .ZN(n8156) );
  AND2_X1 U9416 ( .A1(n9297), .A2(SI_27_), .ZN(n7569) );
  AND2_X1 U9417 ( .A1(n12000), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7570) );
  INV_X1 U9418 ( .A(n8426), .ZN(n7721) );
  NAND2_X1 U9419 ( .A1(n8717), .A2(n8716), .ZN(n12034) );
  INV_X1 U9420 ( .A(n12034), .ZN(n7947) );
  NAND2_X1 U9421 ( .A1(n7835), .A2(n9157), .ZN(n10450) );
  INV_X2 U9422 ( .A(n16567), .ZN(n16570) );
  INV_X1 U9423 ( .A(n10722), .ZN(n8045) );
  INV_X1 U9424 ( .A(n13668), .ZN(n7642) );
  INV_X1 U9425 ( .A(n13632), .ZN(n16366) );
  AND2_X1 U9426 ( .A1(n15385), .A2(n8315), .ZN(n7571) );
  NAND2_X1 U9427 ( .A1(n8816), .A2(n8815), .ZN(n12427) );
  INV_X1 U9428 ( .A(n12427), .ZN(n7955) );
  INV_X1 U9429 ( .A(n16434), .ZN(n7857) );
  NAND2_X1 U9430 ( .A1(n11503), .A2(n13607), .ZN(n8332) );
  INV_X1 U9431 ( .A(n15412), .ZN(n7670) );
  NAND2_X1 U9432 ( .A1(n9870), .A2(n9525), .ZN(n9881) );
  OAI22_X2 U9433 ( .A1(n9789), .A2(n9515), .B1(P1_DATAO_REG_14__SCAN_IN), .B2(
        n10601), .ZN(n9804) );
  INV_X1 U9434 ( .A(n9682), .ZN(n7577) );
  NAND2_X1 U9435 ( .A1(n12779), .A2(n12901), .ZN(n7575) );
  NAND2_X1 U9436 ( .A1(n8149), .A2(n7534), .ZN(n9948) );
  INV_X1 U9437 ( .A(n13400), .ZN(n7627) );
  INV_X1 U9438 ( .A(n9536), .ZN(n8151) );
  NAND2_X1 U9439 ( .A1(n9483), .A2(n9482), .ZN(n9613) );
  OAI21_X1 U9440 ( .B1(n9537), .B2(n9536), .A(n8148), .ZN(n9935) );
  NAND2_X1 U9441 ( .A1(n13781), .A2(n10030), .ZN(n13766) );
  NAND2_X1 U9442 ( .A1(n8003), .A2(n8001), .ZN(n12243) );
  NAND2_X1 U9443 ( .A1(n10010), .A2(n7491), .ZN(n8011) );
  INV_X1 U9444 ( .A(n12300), .ZN(n10006) );
  INV_X2 U9445 ( .A(n9646), .ZN(n13485) );
  AOI21_X1 U9446 ( .B1(n16578), .B2(n13723), .A(n13724), .ZN(n10104) );
  AND2_X2 U9447 ( .A1(n12810), .A2(n12809), .ZN(n12925) );
  NAND2_X1 U9448 ( .A1(n13732), .A2(n13743), .ZN(n13731) );
  NAND2_X1 U9449 ( .A1(n7605), .A2(n12766), .ZN(n13781) );
  NAND2_X1 U9450 ( .A1(n9772), .A2(n12844), .ZN(n13944) );
  INV_X1 U9451 ( .A(n13849), .ZN(n7580) );
  AOI21_X2 U9452 ( .B1(n13742), .B2(n12899), .A(n9989), .ZN(n12734) );
  AOI21_X1 U9453 ( .B1(n12956), .B2(n7479), .A(n12763), .ZN(n12958) );
  NAND2_X1 U9454 ( .A1(n7582), .A2(n7581), .ZN(n13838) );
  NOR2_X1 U9455 ( .A1(n9551), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n7989) );
  NAND2_X1 U9456 ( .A1(n12238), .A2(n12932), .ZN(n12240) );
  NAND2_X1 U9457 ( .A1(n12734), .A2(n12904), .ZN(n12956) );
  NAND2_X1 U9458 ( .A1(n9852), .A2(n12872), .ZN(n13874) );
  INV_X1 U9459 ( .A(n13836), .ZN(n7582) );
  NAND2_X1 U9460 ( .A1(n7957), .A2(n12795), .ZN(n11649) );
  INV_X1 U9461 ( .A(n11651), .ZN(n7957) );
  OAI211_X1 U9462 ( .C1(n7834), .C2(n7833), .A(n7832), .B(n7831), .ZN(n9187)
         );
  OAI22_X1 U9463 ( .A1(n10622), .A2(n14202), .B1(n16420), .B2(n14735), .ZN(
        n10605) );
  OAI22_X2 U9464 ( .A1(n14929), .A2(n12705), .B1(n15048), .B2(n14912), .ZN(
        n14919) );
  NAND2_X1 U9465 ( .A1(n12377), .A2(n12376), .ZN(n12558) );
  OAI21_X1 U9466 ( .B1(n14851), .B2(n8135), .A(n8132), .ZN(n14818) );
  NOR2_X1 U9467 ( .A1(n11452), .A2(n7570), .ZN(n11483) );
  NAND2_X1 U9468 ( .A1(n10761), .A2(n10760), .ZN(n10783) );
  NAND2_X1 U9469 ( .A1(n7652), .A2(n8106), .ZN(n11471) );
  NAND2_X1 U9470 ( .A1(n12174), .A2(n7555), .ZN(n12355) );
  OAI21_X1 U9471 ( .B1(n8102), .B2(n15343), .A(n8096), .ZN(n15227) );
  NAND2_X1 U9472 ( .A1(n10117), .A2(n10116), .ZN(n10357) );
  NAND3_X1 U9473 ( .A1(n8081), .A2(n10526), .A3(n10525), .ZN(n10765) );
  NAND2_X1 U9474 ( .A1(n7586), .A2(n7585), .ZN(n8417) );
  NAND2_X1 U9475 ( .A1(n9240), .A2(n9239), .ZN(n7585) );
  NAND2_X2 U9476 ( .A1(n7522), .A2(n7835), .ZN(n9159) );
  AND2_X1 U9477 ( .A1(n9155), .A2(n9154), .ZN(n7835) );
  NAND2_X1 U9478 ( .A1(n7775), .A2(n8438), .ZN(n8588) );
  NAND2_X1 U9479 ( .A1(n7778), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7633) );
  NAND2_X1 U9480 ( .A1(n8590), .A2(n8438), .ZN(n8614) );
  OAI22_X1 U9481 ( .A1(n9390), .A2(n9391), .B1(n9382), .B2(n9381), .ZN(n7591)
         );
  NAND2_X1 U9482 ( .A1(n7738), .A2(n7533), .ZN(n8672) );
  NAND2_X1 U9483 ( .A1(n8789), .A2(n8788), .ZN(n8474) );
  NAND2_X1 U9484 ( .A1(n9048), .A2(n8261), .ZN(n8259) );
  NAND2_X1 U9485 ( .A1(n8481), .A2(n8482), .ZN(n8868) );
  NAND2_X1 U9486 ( .A1(n7917), .A2(n7923), .ZN(n7916) );
  NAND2_X1 U9487 ( .A1(n7796), .A2(n7442), .ZN(n8484) );
  AND3_X2 U9488 ( .A1(n8871), .A2(n7458), .A3(n7438), .ZN(n15105) );
  NAND2_X1 U9489 ( .A1(n7612), .A2(n7611), .ZN(n7842) );
  OAI21_X1 U9490 ( .B1(n9173), .B2(n9172), .A(n7593), .ZN(n9178) );
  NAND2_X1 U9491 ( .A1(n7595), .A2(n7594), .ZN(n7593) );
  NAND2_X1 U9492 ( .A1(n9173), .A2(n9172), .ZN(n7595) );
  INV_X1 U9493 ( .A(n9179), .ZN(n8388) );
  AOI21_X1 U9494 ( .B1(n9290), .B2(n9289), .A(n7841), .ZN(n7843) );
  NAND2_X1 U9495 ( .A1(n8411), .A2(n8413), .ZN(n9258) );
  INV_X1 U9496 ( .A(n9189), .ZN(n7625) );
  NAND2_X1 U9497 ( .A1(n8525), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n8526) );
  NOR2_X4 U9498 ( .A1(n15847), .A2(n15632), .ZN(n15635) );
  NOR2_X2 U9499 ( .A1(n11981), .A2(n13090), .ZN(n12005) );
  NAND2_X1 U9500 ( .A1(n7934), .A2(n7933), .ZN(P1_U3557) );
  OAI21_X1 U9501 ( .B1(n15834), .B2(n16435), .A(n15833), .ZN(n7882) );
  NAND2_X1 U9502 ( .A1(n8599), .A2(n14208), .ZN(n10711) );
  NAND2_X2 U9503 ( .A1(n8031), .A2(n9157), .ZN(n14884) );
  NAND2_X1 U9504 ( .A1(n8415), .A2(n8416), .ZN(n8541) );
  NAND2_X1 U9505 ( .A1(n10861), .A2(n10862), .ZN(n10872) );
  INV_X1 U9506 ( .A(n15384), .ZN(n7600) );
  NAND2_X1 U9507 ( .A1(n10867), .A2(n7861), .ZN(n7864) );
  INV_X1 U9508 ( .A(n13778), .ZN(n7605) );
  OAI21_X2 U9509 ( .B1(n10049), .B2(n13878), .A(n10048), .ZN(n13724) );
  INV_X1 U9510 ( .A(n16444), .ZN(n13484) );
  NAND2_X2 U9511 ( .A1(n8050), .A2(n8591), .ZN(n16420) );
  INV_X1 U9512 ( .A(n14812), .ZN(n14813) );
  NOR2_X2 U9513 ( .A1(n14955), .A2(n15048), .ZN(n14933) );
  NOR2_X2 U9514 ( .A1(n10987), .A2(n11802), .ZN(n11927) );
  NOR2_X1 U9515 ( .A1(n10716), .A2(n10620), .ZN(n10608) );
  INV_X1 U9516 ( .A(n8176), .ZN(n9758) );
  NAND3_X1 U9517 ( .A1(n8365), .A2(n9458), .A3(n8364), .ZN(n9763) );
  NAND2_X1 U9518 ( .A1(n12107), .A2(n10000), .ZN(n8003) );
  NAND2_X1 U9519 ( .A1(n12805), .A2(n12800), .ZN(n11630) );
  NAND2_X1 U9520 ( .A1(n7606), .A2(n12964), .ZN(P3_U3296) );
  OAI21_X1 U9521 ( .B1(n12959), .B2(n8432), .A(n10745), .ZN(n7606) );
  OAI21_X2 U9522 ( .B1(n8666), .B2(n8046), .A(n8044), .ZN(n10855) );
  AND2_X2 U9523 ( .A1(n8504), .A2(n8503), .ZN(n8871) );
  AOI21_X2 U9524 ( .B1(n14828), .B2(n16507), .A(n7608), .ZN(n15013) );
  INV_X4 U9525 ( .A(n7778), .ZN(n8511) );
  NAND3_X1 U9526 ( .A1(n7742), .A2(n8442), .A3(n7610), .ZN(n7738) );
  NAND2_X1 U9527 ( .A1(n15756), .A2(n15757), .ZN(n8190) );
  NAND3_X1 U9528 ( .A1(n7685), .A2(n10249), .A3(n10166), .ZN(n10123) );
  NAND2_X2 U9529 ( .A1(n11562), .A2(n8184), .ZN(n11583) );
  NAND2_X2 U9530 ( .A1(n8193), .A2(n8191), .ZN(n15866) );
  NOR2_X1 U9531 ( .A1(n9188), .A2(n7854), .ZN(n7626) );
  NAND2_X1 U9532 ( .A1(n7624), .A2(n7852), .ZN(n9200) );
  NAND2_X4 U9533 ( .A1(n12732), .A2(n10036), .ZN(n10928) );
  AND2_X2 U9534 ( .A1(n8346), .A2(n9552), .ZN(n8345) );
  NAND2_X1 U9535 ( .A1(n8347), .A2(n7621), .ZN(n7620) );
  NAND2_X1 U9536 ( .A1(n8403), .A2(n8400), .ZN(n8398) );
  OAI21_X1 U9537 ( .B1(n8269), .B2(n8266), .A(n9402), .ZN(n9442) );
  NAND2_X1 U9538 ( .A1(n7625), .A2(n7626), .ZN(n7624) );
  NAND2_X1 U9539 ( .A1(n7824), .A2(n7823), .ZN(n9173) );
  NAND2_X1 U9540 ( .A1(n7826), .A2(n7827), .ZN(n7823) );
  AND2_X2 U9541 ( .A1(n7647), .A2(n8347), .ZN(n9555) );
  AOI21_X1 U9542 ( .B1(n7618), .B2(n13712), .A(n13711), .ZN(n13713) );
  XNOR2_X1 U9543 ( .A(n13696), .B(n13695), .ZN(n7618) );
  NAND2_X1 U9544 ( .A1(n8011), .A2(n8010), .ZN(n13929) );
  NAND2_X1 U9545 ( .A1(n10014), .A2(n12940), .ZN(n13919) );
  NAND2_X1 U9546 ( .A1(n7993), .A2(n7990), .ZN(n13778) );
  XOR2_X1 U9547 ( .A(n13633), .B(n16366), .Z(n16362) );
  AOI21_X1 U9548 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n13649), .A(n13648), .ZN(
        n13678) );
  INV_X1 U9549 ( .A(n9763), .ZN(n9460) );
  NAND2_X1 U9550 ( .A1(n8527), .A2(n8526), .ZN(n9155) );
  NAND3_X1 U9551 ( .A1(n8388), .A2(n8387), .A3(n7467), .ZN(n7832) );
  INV_X2 U9552 ( .A(n9399), .ZN(n9361) );
  MUX2_X2 U9553 ( .A(n12912), .B(n12911), .S(n12910), .Z(n12917) );
  AOI21_X2 U9554 ( .B1(n12900), .B2(n7470), .A(n7628), .ZN(n12909) );
  OAI21_X1 U9555 ( .B1(n9744), .B2(n9510), .A(n9512), .ZN(n8176) );
  NAND2_X1 U9556 ( .A1(n9490), .A2(n9489), .ZN(n9638) );
  NAND2_X1 U9557 ( .A1(n8175), .A2(n12921), .ZN(n8173) );
  NAND2_X1 U9558 ( .A1(n9537), .A2(n8150), .ZN(n8149) );
  NAND2_X1 U9559 ( .A1(n9493), .A2(n9492), .ZN(n9656) );
  NAND2_X1 U9560 ( .A1(n9497), .A2(n9496), .ZN(n9670) );
  NAND2_X1 U9561 ( .A1(n9869), .A2(n9871), .ZN(n9870) );
  NAND2_X1 U9562 ( .A1(n8047), .A2(n8045), .ZN(n7629) );
  OAI21_X2 U9563 ( .B1(n11157), .B2(n11153), .A(n11154), .ZN(n11377) );
  NAND2_X1 U9564 ( .A1(n9044), .A2(n14638), .ZN(n14693) );
  NAND2_X1 U9565 ( .A1(n8029), .A2(n8028), .ZN(n14618) );
  INV_X1 U9566 ( .A(n8670), .ZN(n8048) );
  NAND2_X1 U9567 ( .A1(n14659), .A2(n8933), .ZN(n14617) );
  NAND2_X1 U9568 ( .A1(n7739), .A2(n8445), .ZN(n8651) );
  MUX2_X1 U9569 ( .A(n9481), .B(n9592), .S(n7778), .Z(n8436) );
  NAND2_X2 U9570 ( .A1(n8245), .A2(n8244), .ZN(n7778) );
  NAND2_X1 U9571 ( .A1(n16304), .A2(n16305), .ZN(n16306) );
  OAI21_X1 U9572 ( .B1(P1_ADDR_REG_1__SCAN_IN), .B2(n16174), .A(n16173), .ZN(
        n16183) );
  NAND2_X1 U9573 ( .A1(n16174), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n7891) );
  INV_X1 U9574 ( .A(n16274), .ZN(n16278) );
  OAI21_X1 U9575 ( .B1(n16220), .B2(n16219), .A(n7895), .ZN(n7894) );
  INV_X1 U9576 ( .A(n8588), .ZN(n8437) );
  NAND2_X1 U9577 ( .A1(n14660), .A2(n8030), .ZN(n14659) );
  INV_X1 U9578 ( .A(n14617), .ZN(n8029) );
  XNOR2_X1 U9579 ( .A(n10938), .B(n11277), .ZN(n11269) );
  AOI22_X1 U9580 ( .A1(n11386), .A2(P3_REG2_REG_7__SCAN_IN), .B1(n11384), .B2(
        n11385), .ZN(n11387) );
  XNOR2_X1 U9581 ( .A(n11383), .B(n11385), .ZN(n11386) );
  AOI21_X1 U9582 ( .B1(n7638), .B2(n7637), .A(n16382), .ZN(n13655) );
  NAND2_X1 U9583 ( .A1(n13650), .A2(n13651), .ZN(n7637) );
  OAI21_X2 U9584 ( .B1(n11397), .B2(n11396), .A(n11395), .ZN(n11681) );
  NAND3_X1 U9585 ( .A1(n7649), .A2(n7542), .A3(n7648), .ZN(n8301) );
  OR2_X1 U9586 ( .A1(n7651), .A2(n13104), .ZN(n7648) );
  NAND2_X1 U9587 ( .A1(n7650), .A2(n13103), .ZN(n7649) );
  NAND2_X1 U9588 ( .A1(n7651), .A2(n13104), .ZN(n7650) );
  NAND2_X1 U9589 ( .A1(n8298), .A2(n8297), .ZN(n7651) );
  NAND2_X2 U9590 ( .A1(n7652), .A2(n7455), .ZN(n10132) );
  NAND2_X1 U9591 ( .A1(n7656), .A2(n7655), .ZN(n8295) );
  INV_X2 U9592 ( .A(n13204), .ZN(n13154) );
  INV_X2 U9593 ( .A(n13290), .ZN(n13155) );
  NAND2_X2 U9594 ( .A1(n10517), .A2(n7668), .ZN(n11173) );
  NAND3_X1 U9595 ( .A1(n13273), .A2(n13272), .A3(n7673), .ZN(n7672) );
  NAND3_X1 U9596 ( .A1(n13229), .A2(n13228), .A3(n7675), .ZN(n7674) );
  NAND2_X1 U9597 ( .A1(n7674), .A2(n7537), .ZN(n8312) );
  NAND2_X1 U9598 ( .A1(n13240), .A2(n13242), .ZN(n7676) );
  NAND2_X1 U9599 ( .A1(n8321), .A2(n7679), .ZN(n7678) );
  NAND2_X1 U9600 ( .A1(n7678), .A2(n7538), .ZN(n8308) );
  NAND2_X1 U9601 ( .A1(n15234), .A2(n7482), .ZN(n7688) );
  NAND2_X1 U9602 ( .A1(n15234), .A2(n7692), .ZN(n7689) );
  AOI21_X1 U9603 ( .B1(n15234), .B2(n15235), .A(n7686), .ZN(n15302) );
  NAND2_X1 U9604 ( .A1(n12055), .A2(n7703), .ZN(n12174) );
  INV_X2 U9605 ( .A(n15136), .ZN(n15255) );
  NAND2_X1 U9606 ( .A1(n15383), .A2(n15252), .ZN(n10498) );
  NOR2_X2 U9607 ( .A1(n15136), .A2(n15793), .ZN(n15252) );
  XNOR2_X2 U9608 ( .A(n7704), .B(n9463), .ZN(n13694) );
  NAND2_X1 U9609 ( .A1(n13526), .A2(n13497), .ZN(n7708) );
  OAI21_X2 U9610 ( .B1(n7709), .B2(n7708), .A(n7706), .ZN(n13500) );
  NAND2_X1 U9611 ( .A1(n12457), .A2(n7714), .ZN(n7712) );
  NAND2_X1 U9612 ( .A1(n7712), .A2(n7531), .ZN(n13374) );
  NAND2_X1 U9613 ( .A1(n7735), .A2(n7734), .ZN(n11093) );
  NAND2_X1 U9614 ( .A1(n7619), .A2(n16428), .ZN(n7734) );
  NAND2_X1 U9615 ( .A1(n11092), .A2(n11093), .ZN(n11091) );
  NAND2_X1 U9616 ( .A1(n11091), .A2(n10948), .ZN(n10950) );
  NOR2_X4 U9617 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n9615) );
  NAND3_X1 U9618 ( .A1(n7742), .A2(n8443), .A3(n8442), .ZN(n7739) );
  NAND2_X1 U9619 ( .A1(n14881), .A2(n7440), .ZN(n7746) );
  NAND2_X1 U9620 ( .A1(n14881), .A2(n14891), .ZN(n12686) );
  NAND2_X1 U9621 ( .A1(n7778), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7754) );
  NAND3_X1 U9622 ( .A1(n7755), .A2(n7754), .A3(n7753), .ZN(n7752) );
  NAND2_X1 U9623 ( .A1(n12641), .A2(n7450), .ZN(n7759) );
  NAND2_X1 U9624 ( .A1(n7759), .A2(n7760), .ZN(n14964) );
  NAND2_X1 U9625 ( .A1(n12192), .A2(n7766), .ZN(n7763) );
  NAND2_X1 U9626 ( .A1(n7763), .A2(n7764), .ZN(n12371) );
  OAI21_X2 U9627 ( .B1(n10892), .B2(n9321), .A(n8676), .ZN(n11934) );
  NAND3_X1 U9628 ( .A1(n15547), .A2(n15569), .A3(n15767), .ZN(n15749) );
  NAND2_X1 U9629 ( .A1(n7777), .A2(n7776), .ZN(n7775) );
  INV_X1 U9630 ( .A(n8229), .ZN(n7780) );
  NAND2_X1 U9631 ( .A1(n7783), .A2(n7782), .ZN(n15861) );
  NAND2_X1 U9632 ( .A1(n7445), .A2(n8229), .ZN(n7783) );
  NAND2_X1 U9633 ( .A1(n7780), .A2(n7782), .ZN(n7779) );
  INV_X1 U9634 ( .A(n7782), .ZN(n7781) );
  NAND2_X1 U9635 ( .A1(n8713), .A2(n7789), .ZN(n7786) );
  OAI21_X1 U9636 ( .B1(n8868), .B2(n8867), .A(n7800), .ZN(n7796) );
  NAND2_X1 U9637 ( .A1(n8870), .A2(n8482), .ZN(n8888) );
  INV_X1 U9638 ( .A(n7795), .ZN(n7794) );
  OAI21_X1 U9639 ( .B1(n15651), .B2(n7815), .A(n7812), .ZN(n15597) );
  NAND2_X1 U9640 ( .A1(n15651), .A2(n7812), .ZN(n7809) );
  AOI21_X1 U9641 ( .B1(n7812), .B2(n7815), .A(n7811), .ZN(n7810) );
  NAND2_X1 U9642 ( .A1(n9166), .A2(n9167), .ZN(n7825) );
  NAND2_X1 U9643 ( .A1(n8388), .A2(n7467), .ZN(n7834) );
  INV_X1 U9644 ( .A(n7836), .ZN(n8411) );
  AOI21_X1 U9645 ( .B1(n8417), .B2(n7837), .A(n7536), .ZN(n7836) );
  NAND2_X1 U9646 ( .A1(n7843), .A2(n7842), .ZN(n7844) );
  NAND2_X1 U9647 ( .A1(n7844), .A2(n7845), .ZN(n8269) );
  INV_X1 U9648 ( .A(n9292), .ZN(n7851) );
  OAI22_X1 U9649 ( .A1(n13290), .A2(n10493), .B1(n13204), .B2(n15404), .ZN(
        n7859) );
  NAND2_X1 U9650 ( .A1(n13311), .A2(n7475), .ZN(n7862) );
  NAND2_X1 U9651 ( .A1(n7864), .A2(n7528), .ZN(n7863) );
  NAND2_X1 U9652 ( .A1(n11203), .A2(n13315), .ZN(n11202) );
  NAND2_X1 U9653 ( .A1(n15763), .A2(n15764), .ZN(n15546) );
  NAND2_X1 U9654 ( .A1(n15866), .A2(n7876), .ZN(n7878) );
  INV_X1 U9655 ( .A(n7878), .ZN(n15662) );
  NOR2_X1 U9656 ( .A1(n15686), .A2(n15557), .ZN(n7880) );
  NAND2_X1 U9657 ( .A1(n11583), .A2(n7881), .ZN(n11806) );
  INV_X1 U9658 ( .A(n16240), .ZN(n7883) );
  NOR2_X2 U9659 ( .A1(n16333), .A2(n16334), .ZN(n16347) );
  OR2_X1 U9660 ( .A1(n10956), .A2(n10955), .ZN(n7896) );
  NAND2_X1 U9661 ( .A1(n10977), .A2(n7897), .ZN(n10959) );
  AND2_X1 U9662 ( .A1(n7898), .A2(n10958), .ZN(n7897) );
  NAND2_X1 U9663 ( .A1(n10956), .A2(n10955), .ZN(n7898) );
  NAND3_X1 U9664 ( .A1(n7904), .A2(n7907), .A3(n7901), .ZN(n11233) );
  NAND3_X1 U9665 ( .A1(n7904), .A2(n7902), .A3(n7901), .ZN(n11405) );
  INV_X1 U9666 ( .A(n8487), .ZN(n7917) );
  NAND3_X1 U9667 ( .A1(n7921), .A2(n7918), .A3(n7916), .ZN(n8981) );
  AOI21_X2 U9668 ( .B1(n15832), .B2(n16458), .A(n7935), .ZN(n15833) );
  INV_X2 U9669 ( .A(n7937), .ZN(n15651) );
  NAND2_X1 U9670 ( .A1(n8812), .A2(n8271), .ZN(n7941) );
  NAND2_X1 U9671 ( .A1(n7941), .A2(n7942), .ZN(n8480) );
  NAND2_X1 U9672 ( .A1(n7941), .A2(n7940), .ZN(n8482) );
  NAND3_X1 U9673 ( .A1(n7943), .A2(n7944), .A3(n8609), .ZN(n8611) );
  NAND2_X1 U9674 ( .A1(n7943), .A2(n8609), .ZN(n7945) );
  NAND2_X1 U9675 ( .A1(n7946), .A2(n10150), .ZN(n7943) );
  NAND2_X1 U9676 ( .A1(n7945), .A2(n8568), .ZN(n8569) );
  INV_X1 U9677 ( .A(n8614), .ZN(n7946) );
  NAND3_X1 U9678 ( .A1(n16617), .A2(n7954), .A3(n12078), .ZN(n12560) );
  NOR2_X2 U9679 ( .A1(n12651), .A2(n15068), .ZN(n14985) );
  NAND2_X1 U9680 ( .A1(n9607), .A2(n12788), .ZN(n11651) );
  XNOR2_X1 U9681 ( .A(n7958), .B(n12798), .ZN(n12795) );
  OAI21_X1 U9682 ( .B1(n7607), .B2(n7965), .A(n7963), .ZN(n12474) );
  NAND2_X1 U9683 ( .A1(n7961), .A2(n7959), .ZN(n9751) );
  AOI21_X1 U9684 ( .B1(n7963), .B2(n7965), .A(n7960), .ZN(n7959) );
  NAND2_X1 U9685 ( .A1(n12240), .A2(n7963), .ZN(n7961) );
  OAI21_X1 U9686 ( .B1(n7444), .B2(n7965), .A(n12834), .ZN(n7964) );
  NAND2_X1 U9687 ( .A1(n12934), .A2(n12829), .ZN(n7965) );
  NAND2_X1 U9688 ( .A1(n13874), .A2(n7971), .ZN(n7967) );
  NAND2_X1 U9689 ( .A1(n11746), .A2(n7977), .ZN(n7974) );
  NAND2_X1 U9690 ( .A1(n7974), .A2(n7975), .ZN(n12238) );
  NAND3_X1 U9691 ( .A1(n12732), .A2(n13671), .A3(n7619), .ZN(n9617) );
  AND2_X2 U9692 ( .A1(n13919), .A2(n10015), .ZN(n13903) );
  NAND2_X1 U9693 ( .A1(n13822), .A2(n7994), .ZN(n7993) );
  OAI21_X1 U9694 ( .B1(n13822), .B2(n7478), .A(n10027), .ZN(n13804) );
  NAND2_X1 U9695 ( .A1(n8004), .A2(n7532), .ZN(n13965) );
  NAND2_X1 U9696 ( .A1(n10006), .A2(n8005), .ZN(n8004) );
  NAND2_X1 U9697 ( .A1(n13875), .A2(n8015), .ZN(n8014) );
  NAND2_X2 U9698 ( .A1(n8014), .A2(n8012), .ZN(n13853) );
  NAND2_X2 U9699 ( .A1(n10928), .A2(n10165), .ZN(n9644) );
  NAND2_X1 U9700 ( .A1(n14158), .A2(n14157), .ZN(n8021) );
  NAND2_X1 U9701 ( .A1(n14652), .A2(n9018), .ZN(n9044) );
  NAND2_X1 U9702 ( .A1(n8022), .A2(n8024), .ZN(n12609) );
  NAND3_X1 U9703 ( .A1(n12087), .A2(n8826), .A3(n12132), .ZN(n8022) );
  AND2_X1 U9704 ( .A1(n9130), .A2(n8032), .ZN(n11324) );
  OAI21_X1 U9705 ( .B1(n8897), .B2(n8041), .A(n8038), .ZN(n8928) );
  NAND2_X1 U9706 ( .A1(n8871), .A2(n8514), .ZN(n8889) );
  NAND2_X1 U9707 ( .A1(n8871), .A2(n8049), .ZN(n8522) );
  NAND2_X1 U9708 ( .A1(n13851), .A2(n12879), .ZN(n13836) );
  OAI211_X2 U9709 ( .C1(n7430), .C2(n10339), .A(n9597), .B(n9596), .ZN(n11032)
         );
  OAI211_X1 U9710 ( .C1(n8175), .C2(n11534), .A(n8174), .B(n8173), .ZN(n12959)
         );
  XNOR2_X2 U9711 ( .A(n14735), .B(n16420), .ZN(n10622) );
  NAND2_X4 U9712 ( .A1(n8802), .A2(n10165), .ZN(n9357) );
  OAI21_X2 U9713 ( .B1(n12568), .B2(n8053), .A(n7480), .ZN(n12644) );
  INV_X1 U9714 ( .A(n12687), .ZN(n8058) );
  NAND2_X1 U9715 ( .A1(n10816), .A2(n10815), .ZN(n8063) );
  NAND3_X1 U9716 ( .A1(n8059), .A2(n10999), .A3(n8061), .ZN(n11346) );
  NAND2_X1 U9717 ( .A1(n10816), .A2(n8060), .ZN(n8059) );
  NAND2_X1 U9718 ( .A1(n8062), .A2(n10995), .ZN(n8061) );
  NAND3_X1 U9719 ( .A1(n8077), .A2(n8074), .A3(n14981), .ZN(n8073) );
  XNOR2_X2 U9720 ( .A(n8079), .B(n8539), .ZN(n15115) );
  NAND3_X1 U9721 ( .A1(n8871), .A2(n7438), .A3(n8509), .ZN(n8080) );
  AOI21_X1 U9722 ( .B1(n10525), .B2(n10526), .A(n8081), .ZN(n10542) );
  XNOR2_X1 U9723 ( .A(n10752), .B(n10751), .ZN(n8081) );
  OAI21_X1 U9724 ( .B1(n15287), .B2(n8087), .A(n8084), .ZN(n15329) );
  NAND2_X1 U9725 ( .A1(n15280), .A2(n8092), .ZN(n8091) );
  AND2_X1 U9726 ( .A1(n8102), .A2(n8101), .ZN(n15345) );
  NAND2_X1 U9727 ( .A1(n10117), .A2(n8110), .ZN(n10336) );
  NAND2_X1 U9728 ( .A1(n10117), .A2(n8108), .ZN(n8107) );
  INV_X1 U9729 ( .A(n8114), .ZN(n15309) );
  NAND2_X1 U9730 ( .A1(n8115), .A2(n7529), .ZN(n12055) );
  INV_X2 U9731 ( .A(n9357), .ZN(n8910) );
  NAND2_X2 U9732 ( .A1(n8572), .A2(n8116), .ZN(n10716) );
  NAND2_X1 U9733 ( .A1(n12649), .A2(n7527), .ZN(n12698) );
  NAND2_X1 U9734 ( .A1(n11341), .A2(n8122), .ZN(n8119) );
  OAI21_X1 U9735 ( .B1(n14851), .B2(n12713), .A(n12714), .ZN(n14833) );
  OAI21_X1 U9736 ( .B1(n12032), .B2(n8139), .A(n8137), .ZN(n12145) );
  OAI21_X2 U9737 ( .B1(n9822), .B2(n8156), .A(n8152), .ZN(n9869) );
  NAND2_X1 U9738 ( .A1(n9881), .A2(n7559), .ZN(n8171) );
  NAND2_X2 U9739 ( .A1(n9533), .A2(n9532), .ZN(n9917) );
  OR2_X2 U9740 ( .A1(n9712), .A2(n9711), .ZN(n9714) );
  OAI21_X2 U9741 ( .B1(n8177), .B2(n9644), .A(n9951), .ZN(n13996) );
  NAND2_X2 U9742 ( .A1(n11068), .A2(n11067), .ZN(n11562) );
  NAND2_X1 U9743 ( .A1(n11861), .A2(n8186), .ZN(n11958) );
  NAND2_X1 U9744 ( .A1(n15601), .A2(n8198), .ZN(n8194) );
  OAI211_X1 U9745 ( .C1(n15601), .C2(n8201), .A(n8199), .B(n8194), .ZN(n15834)
         );
  OAI21_X1 U9746 ( .B1(n15834), .B2(n8197), .A(n8195), .ZN(P1_U3525) );
  OAI21_X2 U9747 ( .B1(n10872), .B2(n7571), .A(n10862), .ZN(n11137) );
  NOR2_X2 U9748 ( .A1(n11363), .A2(n11362), .ZN(n11366) );
  NAND2_X1 U9749 ( .A1(n15635), .A2(n8207), .ZN(n15584) );
  INV_X1 U9750 ( .A(n15607), .ZN(n15585) );
  NAND2_X1 U9751 ( .A1(n12004), .A2(n8217), .ZN(n8216) );
  NAND2_X1 U9752 ( .A1(n11059), .A2(n8223), .ZN(n8222) );
  NAND2_X1 U9753 ( .A1(n15713), .A2(n8230), .ZN(n8229) );
  NAND2_X1 U9754 ( .A1(n8240), .A2(n8239), .ZN(P1_U3523) );
  OR2_X1 U9755 ( .A1(n16570), .A2(n13013), .ZN(n8239) );
  XNOR2_X1 U9756 ( .A(n15612), .B(n15624), .ZN(n8243) );
  INV_X1 U9757 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n15525) );
  NAND4_X1 U9758 ( .A1(n16349), .A2(n16385), .A3(P1_ADDR_REG_19__SCAN_IN), 
        .A4(P2_ADDR_REG_19__SCAN_IN), .ZN(n8244) );
  NAND4_X1 U9759 ( .A1(n8433), .A2(n8434), .A3(n15525), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n8245) );
  NAND2_X1 U9760 ( .A1(n8246), .A2(n8247), .ZN(n8711) );
  NAND2_X1 U9761 ( .A1(n8672), .A2(n8249), .ZN(n8246) );
  NAND2_X1 U9762 ( .A1(n13203), .A2(n8255), .ZN(n8254) );
  NAND2_X1 U9763 ( .A1(n9048), .A2(n9047), .ZN(n9071) );
  NAND3_X1 U9764 ( .A1(n8267), .A2(n7477), .A3(n9397), .ZN(n8266) );
  OAI21_X1 U9765 ( .B1(n8936), .B2(n8935), .A(n8938), .ZN(n8958) );
  INV_X1 U9766 ( .A(n8284), .ZN(n8283) );
  NAND2_X1 U9767 ( .A1(n8285), .A2(n8957), .ZN(n8284) );
  NAND2_X1 U9768 ( .A1(n13077), .A2(n8286), .ZN(n8291) );
  INV_X1 U9769 ( .A(n13076), .ZN(n8289) );
  INV_X1 U9770 ( .A(n13087), .ZN(n8296) );
  NAND3_X1 U9771 ( .A1(n13098), .A2(n13097), .A3(n7540), .ZN(n8298) );
  INV_X1 U9772 ( .A(n13099), .ZN(n8299) );
  INV_X1 U9773 ( .A(n13106), .ZN(n8302) );
  NAND3_X1 U9774 ( .A1(n13120), .A2(n13119), .A3(n7539), .ZN(n8304) );
  INV_X1 U9775 ( .A(n13132), .ZN(n8305) );
  INV_X1 U9776 ( .A(n13193), .ZN(n8309) );
  INV_X1 U9777 ( .A(n13253), .ZN(n8313) );
  NAND2_X1 U9778 ( .A1(n8316), .A2(n7449), .ZN(n15385) );
  AND2_X1 U9779 ( .A1(n8314), .A2(n10353), .ZN(n8316) );
  NAND2_X1 U9780 ( .A1(n13310), .A2(n15384), .ZN(n13026) );
  NAND3_X1 U9781 ( .A1(n13152), .A2(n13151), .A3(n8318), .ZN(n8321) );
  INV_X1 U9782 ( .A(n13166), .ZN(n8320) );
  NAND3_X1 U9783 ( .A1(n8324), .A2(n8325), .A3(n13276), .ZN(n8322) );
  INV_X1 U9784 ( .A(n10132), .ZN(n8326) );
  NOR2_X1 U9785 ( .A1(n10132), .A2(n8329), .ZN(n10345) );
  NAND2_X1 U9786 ( .A1(n11710), .A2(n11711), .ZN(n12157) );
  OAI211_X1 U9787 ( .C1(n13573), .C2(n8340), .A(n8337), .B(n8335), .ZN(n13435)
         );
  NAND2_X1 U9788 ( .A1(n13573), .A2(n8336), .ZN(n8335) );
  NOR2_X1 U9789 ( .A1(n13429), .A2(n8338), .ZN(n8336) );
  OAI22_X1 U9790 ( .A1(n8339), .A2(n8338), .B1(n13429), .B2(n8341), .ZN(n8337)
         );
  NOR2_X1 U9791 ( .A1(n13429), .A2(n13453), .ZN(n8339) );
  NAND2_X1 U9792 ( .A1(n13453), .A2(n13429), .ZN(n8340) );
  INV_X2 U9793 ( .A(n9765), .ZN(n8347) );
  NAND2_X1 U9794 ( .A1(n13460), .A2(n7526), .ZN(n8348) );
  NAND2_X1 U9795 ( .A1(n13382), .A2(n13934), .ZN(n8363) );
  NAND2_X1 U9796 ( .A1(n8369), .A2(n8370), .ZN(n13404) );
  NAND2_X1 U9797 ( .A1(n13389), .A2(n13388), .ZN(n13491) );
  AND2_X2 U9798 ( .A1(n9555), .A2(n8379), .ZN(n9577) );
  INV_X4 U9799 ( .A(n9159), .ZN(n9371) );
  NAND2_X1 U9800 ( .A1(n14737), .A2(n10660), .ZN(n9421) );
  OAI21_X1 U9801 ( .B1(n14737), .B2(n9159), .A(n8382), .ZN(n8384) );
  INV_X1 U9802 ( .A(n8383), .ZN(n8382) );
  OAI21_X1 U9803 ( .B1(n10660), .B2(n9159), .A(n11319), .ZN(n8383) );
  NAND2_X1 U9804 ( .A1(n8384), .A2(n9158), .ZN(n9163) );
  NOR2_X1 U9805 ( .A1(n9213), .A2(n9212), .ZN(n9214) );
  INV_X1 U9806 ( .A(n9206), .ZN(n8386) );
  INV_X1 U9807 ( .A(n9182), .ZN(n8387) );
  INV_X1 U9808 ( .A(n9283), .ZN(n8401) );
  NAND2_X1 U9809 ( .A1(n9279), .A2(n9280), .ZN(n8403) );
  INV_X1 U9810 ( .A(n8404), .ZN(n9240) );
  OR2_X1 U9811 ( .A1(n12995), .A2(n13373), .ZN(n15805) );
  OR2_X2 U9812 ( .A1(n12145), .A2(n12144), .ZN(n12072) );
  NAND2_X1 U9813 ( .A1(n9932), .A2(n12781), .ZN(n13776) );
  NAND2_X1 U9814 ( .A1(n13790), .A2(n12780), .ZN(n9932) );
  NAND2_X1 U9815 ( .A1(n10873), .A2(n10872), .ZN(n11125) );
  CLKBUF_X1 U9816 ( .A(n13929), .Z(n13952) );
  XNOR2_X2 U9817 ( .A(n10716), .B(n14734), .ZN(n10610) );
  OR2_X1 U9818 ( .A1(n13284), .A2(n16413), .ZN(n10419) );
  CLKBUF_X1 U9819 ( .A(n13440), .Z(n13442) );
  NAND2_X1 U9820 ( .A1(n9575), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9576) );
  XNOR2_X1 U9821 ( .A(n15380), .B(n13053), .ZN(n13311) );
  NAND2_X1 U9822 ( .A1(n9413), .A2(n9412), .ZN(n9454) );
  NAND2_X1 U9823 ( .A1(n9442), .A2(n9411), .ZN(n9412) );
  AND2_X1 U9824 ( .A1(n11524), .A2(n13946), .ZN(n13958) );
  NAND2_X1 U9825 ( .A1(n16587), .A2(n14040), .ZN(n14051) );
  INV_X1 U9826 ( .A(n14051), .ZN(n10089) );
  INV_X1 U9827 ( .A(n13606), .ZN(n11644) );
  NOR2_X1 U9828 ( .A1(n11943), .A2(n12925), .ZN(n8424) );
  INV_X1 U9829 ( .A(n15687), .ZN(n15556) );
  NOR3_X1 U9830 ( .A1(n14886), .A2(n14885), .A3(n14884), .ZN(n8425) );
  INV_X1 U9831 ( .A(n14707), .ZN(n14686) );
  AND2_X2 U9832 ( .A1(n11054), .A2(n11118), .ZN(n16469) );
  INV_X2 U9833 ( .A(n16605), .ZN(n15812) );
  AND2_X1 U9834 ( .A1(n12455), .A2(n13604), .ZN(n8426) );
  NOR2_X1 U9835 ( .A1(n10025), .A2(n10024), .ZN(n8427) );
  OR2_X1 U9836 ( .A1(n13377), .A2(n13376), .ZN(n8429) );
  INV_X1 U9837 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10115) );
  INV_X1 U9838 ( .A(n12934), .ZN(n12306) );
  AND4_X1 U9839 ( .A1(n9125), .A2(n8514), .A3(n8906), .A4(n8515), .ZN(n8430)
         );
  AND3_X1 U9840 ( .A1(n9445), .A2(n9444), .A3(n12727), .ZN(n8431) );
  INV_X1 U9841 ( .A(P1_RD_REG_SCAN_IN), .ZN(n8434) );
  INV_X1 U9842 ( .A(n9341), .ZN(n8836) );
  INV_X1 U9843 ( .A(n13907), .ZN(n10016) );
  INV_X1 U9844 ( .A(n13824), .ZN(n13794) );
  AND3_X1 U9845 ( .A1(n9924), .A2(n9923), .A3(n9922), .ZN(n13824) );
  AND4_X1 U9846 ( .A1(n12958), .A2(n12957), .A3(n12956), .A4(n12955), .ZN(
        n8432) );
  AND2_X1 U9847 ( .A1(n13026), .A2(n13025), .ZN(n13038) );
  AND2_X1 U9848 ( .A1(n13043), .A2(n13042), .ZN(n13039) );
  OAI21_X1 U9849 ( .B1(n9403), .B2(n10660), .A(n9159), .ZN(n9160) );
  INV_X1 U9850 ( .A(n9160), .ZN(n9161) );
  NAND2_X1 U9851 ( .A1(n14737), .A2(n9161), .ZN(n9162) );
  INV_X1 U9852 ( .A(n12947), .ZN(n12897) );
  INV_X1 U9853 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8499) );
  INV_X1 U9854 ( .A(n13949), .ZN(n10012) );
  INV_X1 U9855 ( .A(n8522), .ZN(n8517) );
  OR2_X1 U9856 ( .A1(n9649), .A2(n9586), .ZN(n9587) );
  INV_X1 U9857 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8433) );
  INV_X1 U9858 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n10129) );
  NAND2_X1 U9859 ( .A1(n13605), .A2(n12385), .ZN(n12386) );
  INV_X1 U9860 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n14273) );
  INV_X1 U9861 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n14464) );
  INV_X1 U9862 ( .A(n13750), .ZN(n10033) );
  NOR2_X1 U9863 ( .A1(n13754), .A2(n13970), .ZN(n10046) );
  INV_X1 U9864 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n9459) );
  AND2_X1 U9865 ( .A1(n9006), .A2(n9005), .ZN(n9030) );
  INV_X1 U9866 ( .A(n8914), .ZN(n8537) );
  XNOR2_X1 U9867 ( .A(n10474), .B(n15221), .ZN(n10476) );
  INV_X1 U9868 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11304) );
  INV_X1 U9869 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n11070) );
  INV_X1 U9870 ( .A(n11471), .ZN(n10117) );
  INV_X1 U9871 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n14587) );
  INV_X1 U9872 ( .A(n11904), .ZN(n11893) );
  INV_X1 U9873 ( .A(n9663), .ZN(n9561) );
  INV_X1 U9874 ( .A(n13694), .ZN(n13706) );
  INV_X1 U9875 ( .A(n8967), .ZN(n8965) );
  INV_X1 U9876 ( .A(n8943), .ZN(n8941) );
  AND2_X1 U9877 ( .A1(n9076), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9138) );
  OR2_X1 U9878 ( .A1(n8916), .A2(n8555), .ZN(n8557) );
  NAND2_X1 U9879 ( .A1(n8537), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8916) );
  AND2_X1 U9880 ( .A1(n10269), .A2(n9446), .ZN(n10445) );
  INV_X1 U9881 ( .A(n12520), .ZN(n12517) );
  INV_X1 U9882 ( .A(n13244), .ZN(n13258) );
  INV_X1 U9883 ( .A(n13320), .ZN(n11563) );
  NAND2_X1 U9884 ( .A1(n8464), .A2(SI_10_), .ZN(n8468) );
  INV_X1 U9885 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n14579) );
  INV_X1 U9886 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n16349) );
  NAND2_X1 U9887 ( .A1(n11654), .A2(n11034), .ZN(n11191) );
  INV_X1 U9888 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n11254) );
  INV_X1 U9889 ( .A(n13920), .ZN(n13594) );
  INV_X1 U9890 ( .A(n16036), .ZN(n16364) );
  AND4_X1 U9891 ( .A1(n9892), .A2(n9891), .A3(n9890), .A4(n9889), .ZN(n13867)
         );
  INV_X1 U9892 ( .A(n13890), .ZN(n13887) );
  INV_X1 U9893 ( .A(n12940), .ZN(n13917) );
  AND2_X1 U9894 ( .A1(n10096), .A2(n12763), .ZN(n13878) );
  AND2_X1 U9895 ( .A1(n13706), .A2(n11281), .ZN(n12920) );
  OR2_X1 U9896 ( .A1(n8837), .A2(n12129), .ZN(n8858) );
  NAND2_X1 U9897 ( .A1(n8965), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n9004) );
  INV_X1 U9898 ( .A(n14718), .ZN(n14177) );
  NAND2_X1 U9899 ( .A1(n8941), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8967) );
  CLKBUF_X3 U9900 ( .A(n8598), .Z(n9075) );
  OR2_X1 U9901 ( .A1(n9148), .A2(n9446), .ZN(n14650) );
  AND2_X1 U9902 ( .A1(n9133), .A2(n16040), .ZN(n9129) );
  INV_X1 U9903 ( .A(n9406), .ZN(n9407) );
  OR2_X1 U9904 ( .A1(n14643), .A2(n9341), .ZN(n9039) );
  OR2_X1 U9905 ( .A1(n8892), .A2(n12534), .ZN(n8914) );
  INV_X1 U9906 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10368) );
  OR2_X1 U9907 ( .A1(n16123), .A2(n16122), .ZN(n16125) );
  INV_X1 U9908 ( .A(n9155), .ZN(n9441) );
  INV_X1 U9909 ( .A(n15062), .ZN(n14995) );
  INV_X1 U9910 ( .A(n14722), .ZN(n12571) );
  AND2_X1 U9911 ( .A1(n9130), .A2(n9446), .ZN(n15079) );
  AND2_X1 U9912 ( .A1(n10458), .A2(n10457), .ZN(n14949) );
  INV_X1 U9913 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n15106) );
  INV_X1 U9914 ( .A(n11619), .ZN(n11620) );
  OR2_X1 U9915 ( .A1(n10423), .A2(n10416), .ZN(n15264) );
  NAND2_X1 U9916 ( .A1(n15997), .A2(n12984), .ZN(n12995) );
  AND2_X1 U9917 ( .A1(n13196), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n13209) );
  AND2_X1 U9918 ( .A1(n13138), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13158) );
  OR2_X1 U9919 ( .A1(n12413), .A2(n12412), .ZN(n13122) );
  INV_X1 U9920 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n16192) );
  OR2_X1 U9921 ( .A1(n12334), .A2(n12333), .ZN(n12335) );
  INV_X1 U9922 ( .A(n15830), .ZN(n13305) );
  INV_X1 U9923 ( .A(n15741), .ZN(n15549) );
  INV_X1 U9924 ( .A(n15910), .ZN(n15915) );
  OR2_X1 U9925 ( .A1(n16493), .A2(n12984), .ZN(n10859) );
  INV_X1 U9926 ( .A(n12980), .ZN(n10409) );
  INV_X1 U9927 ( .A(n16556), .ZN(n16490) );
  OR2_X1 U9928 ( .A1(n12995), .A2(n10417), .ZN(n16389) );
  XNOR2_X1 U9929 ( .A(n8479), .B(SI_15_), .ZN(n8849) );
  OAI21_X1 U9930 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n16310), .A(n16309), .ZN(
        n16314) );
  INV_X1 U9931 ( .A(n13593), .ZN(n13566) );
  INV_X1 U9932 ( .A(n13448), .ZN(n13590) );
  AND2_X1 U9933 ( .A1(n12743), .A2(n12742), .ZN(n13717) );
  INV_X1 U9934 ( .A(n13867), .ZN(n13834) );
  INV_X1 U9935 ( .A(n16382), .ZN(n13712) );
  AND2_X1 U9936 ( .A1(n11037), .A2(n12910), .ZN(n13967) );
  INV_X1 U9937 ( .A(n12814), .ZN(n12164) );
  INV_X1 U9938 ( .A(n13946), .ZN(n13980) );
  AND2_X1 U9939 ( .A1(n10081), .A2(n10080), .ZN(n11517) );
  INV_X1 U9940 ( .A(n14139), .ZN(n10106) );
  AND2_X1 U9941 ( .A1(n13976), .A2(n13975), .ZN(n14132) );
  INV_X1 U9942 ( .A(n14109), .ZN(n14134) );
  OR2_X1 U9943 ( .A1(n14052), .A2(n16485), .ZN(n16578) );
  XNOR2_X1 U9944 ( .A(n10075), .B(n10076), .ZN(n10926) );
  AND2_X1 U9945 ( .A1(n9525), .A2(n9524), .ZN(n9871) );
  INV_X1 U9946 ( .A(n9826), .ZN(n9840) );
  AND2_X1 U9947 ( .A1(n9129), .A2(n9127), .ZN(n14707) );
  OR2_X1 U9948 ( .A1(n14194), .A2(n9341), .ZN(n9147) );
  NAND2_X1 U9949 ( .A1(n8894), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8582) );
  OR2_X1 U9950 ( .A1(n16087), .A2(P2_U3088), .ZN(n16127) );
  INV_X1 U9951 ( .A(n11858), .ZN(n16148) );
  INV_X1 U9952 ( .A(n16114), .ZN(n16152) );
  NAND2_X1 U9953 ( .A1(n12694), .A2(n12693), .ZN(n12695) );
  INV_X1 U9954 ( .A(n12688), .ZN(n14859) );
  INV_X1 U9955 ( .A(n16511), .ZN(n14922) );
  AND2_X1 U9956 ( .A1(n12375), .A2(n12264), .ZN(n12425) );
  INV_X1 U9957 ( .A(n14829), .ZN(n16519) );
  INV_X1 U9958 ( .A(n14926), .ZN(n16508) );
  INV_X1 U9959 ( .A(n14949), .ZN(n14981) );
  INV_X1 U9960 ( .A(n15079), .ZN(n16616) );
  INV_X1 U9961 ( .A(n16621), .ZN(n15082) );
  OR2_X1 U9962 ( .A1(n16507), .A2(n16610), .ZN(n16621) );
  AND3_X1 U9963 ( .A1(n11318), .A2(n16032), .A3(n10447), .ZN(n10603) );
  AND2_X1 U9964 ( .A1(n10273), .A2(n9414), .ZN(n10270) );
  INV_X1 U9965 ( .A(n15398), .ZN(n15517) );
  INV_X1 U9966 ( .A(n15511), .ZN(n15477) );
  INV_X1 U9967 ( .A(n15512), .ZN(n15516) );
  AND2_X1 U9968 ( .A1(n16386), .A2(n12993), .ZN(n15910) );
  INV_X1 U9969 ( .A(n15542), .ZN(n15816) );
  XNOR2_X1 U9970 ( .A(n11173), .B(n15382), .ZN(n13312) );
  OR2_X1 U9971 ( .A1(n10424), .A2(n10859), .ZN(n16395) );
  AND2_X1 U9972 ( .A1(n16454), .A2(n16493), .ZN(n16435) );
  INV_X1 U9973 ( .A(n16458), .ZN(n16558) );
  INV_X1 U9974 ( .A(n16435), .ZN(n16564) );
  NAND2_X1 U9975 ( .A1(n10880), .A2(n10879), .ZN(n16458) );
  NOR2_X1 U9976 ( .A1(n10182), .A2(n15985), .ZN(n10401) );
  XNOR2_X1 U9977 ( .A(n9295), .B(n9072), .ZN(n15118) );
  INV_X1 U9978 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n16167) );
  AND2_X1 U9979 ( .A1(n10963), .A2(n10962), .ZN(n16036) );
  AND2_X1 U9980 ( .A1(n10748), .A2(n10747), .ZN(n13448) );
  INV_X1 U9981 ( .A(n13596), .ZN(n13582) );
  AND2_X1 U9982 ( .A1(n12743), .A2(n10044), .ZN(n12913) );
  OAI211_X1 U9983 ( .C1(n7436), .C2(n13821), .A(n9914), .B(n9913), .ZN(n13833)
         );
  INV_X1 U9984 ( .A(n13550), .ZN(n13955) );
  INV_X1 U9985 ( .A(P3_U3897), .ZN(n13606) );
  INV_X1 U9986 ( .A(n13707), .ZN(n16367) );
  AND2_X1 U9987 ( .A1(n13737), .A2(n13736), .ZN(n13990) );
  NAND2_X1 U9988 ( .A1(n13977), .A2(n11538), .ZN(n13963) );
  NAND2_X1 U9989 ( .A1(n13977), .A2(n11635), .ZN(n13984) );
  NAND2_X1 U9990 ( .A1(n10088), .A2(n10089), .ZN(n10090) );
  INV_X1 U9991 ( .A(n16587), .ZN(n16585) );
  AND3_X2 U9992 ( .A1(n10086), .A2(n11517), .A3(n10085), .ZN(n16587) );
  NAND2_X1 U9993 ( .A1(n16590), .A2(n14040), .ZN(n14139) );
  INV_X1 U9994 ( .A(n16590), .ZN(n16588) );
  AND2_X1 U9995 ( .A1(n10061), .A2(n10060), .ZN(n14141) );
  AND2_X1 U9996 ( .A1(n10926), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14140) );
  INV_X1 U9997 ( .A(SI_16_), .ZN(n14429) );
  INV_X1 U9998 ( .A(SI_12_), .ZN(n14236) );
  INV_X1 U9999 ( .A(n14691), .ZN(n14705) );
  NAND2_X1 U10000 ( .A1(n9147), .A2(n9146), .ZN(n14839) );
  NAND2_X1 U10001 ( .A1(n8991), .A2(n8990), .ZN(n14914) );
  OR2_X1 U10002 ( .A1(n8862), .A2(n8861), .ZN(n14721) );
  OR2_X1 U10003 ( .A1(n10307), .A2(n15119), .ZN(n16114) );
  OR2_X1 U10004 ( .A1(n10307), .A2(n10306), .ZN(n11858) );
  OR2_X1 U10005 ( .A1(n11787), .A2(n11851), .ZN(n14926) );
  AND2_X1 U10006 ( .A1(n12647), .A2(n12646), .ZN(n15070) );
  AND2_X1 U10007 ( .A1(n14829), .A2(n11796), .ZN(n14892) );
  OR2_X1 U10008 ( .A1(n16522), .A2(n11320), .ZN(n14829) );
  NAND2_X1 U10009 ( .A1(n10603), .A2(n16039), .ZN(n16623) );
  OR2_X1 U10010 ( .A1(n16037), .A2(n16034), .ZN(n16035) );
  NAND2_X1 U10011 ( .A1(n9118), .A2(n9117), .ZN(n16039) );
  XNOR2_X1 U10012 ( .A(n9112), .B(n9111), .ZN(n15130) );
  INV_X1 U10013 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11495) );
  INV_X1 U10014 ( .A(n12470), .ZN(n15131) );
  INV_X1 U10015 ( .A(n15365), .ZN(n15340) );
  OR2_X1 U10016 ( .A1(n10423), .A2(n10408), .ZN(n15367) );
  INV_X1 U10017 ( .A(n15636), .ZN(n15370) );
  OR2_X1 U10018 ( .A1(n16164), .A2(n16159), .ZN(n15398) );
  INV_X1 U10019 ( .A(n16162), .ZN(n15524) );
  INV_X1 U10020 ( .A(n15711), .ZN(n15821) );
  OR3_X1 U10021 ( .A1(n15908), .A2(n15907), .A3(n15906), .ZN(n15962) );
  NAND2_X1 U10022 ( .A1(n11054), .A2(n11053), .ZN(n16567) );
  INV_X2 U10023 ( .A(n16000), .ZN(n16031) );
  INV_X1 U10024 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11012) );
  AND2_X1 U10025 ( .A1(n14140), .A2(n10141), .ZN(P3_U3897) );
  NAND2_X1 U10026 ( .A1(n8435), .A2(SI_1_), .ZN(n8438) );
  INV_X1 U10027 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9592) );
  INV_X2 U10028 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9481) );
  INV_X1 U10029 ( .A(SI_0_), .ZN(n10339) );
  NOR2_X1 U10030 ( .A1(n8436), .A2(n10339), .ZN(n8586) );
  NAND2_X1 U10031 ( .A1(n8437), .A2(n8586), .ZN(n8590) );
  INV_X1 U10032 ( .A(SI_2_), .ZN(n10150) );
  NOR2_X1 U10033 ( .A1(n8568), .A2(n10150), .ZN(n8613) );
  INV_X1 U10034 ( .A(n8613), .ZN(n8439) );
  NAND2_X1 U10035 ( .A1(n8439), .A2(n8629), .ZN(n8444) );
  INV_X1 U10036 ( .A(n8612), .ZN(n8440) );
  NAND2_X1 U10037 ( .A1(n8440), .A2(n8629), .ZN(n8443) );
  MUX2_X1 U10038 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8511), .Z(n8441) );
  NAND2_X1 U10039 ( .A1(n8441), .A2(SI_4_), .ZN(n8445) );
  OAI21_X1 U10040 ( .B1(n8441), .B2(SI_4_), .A(n8445), .ZN(n8631) );
  MUX2_X1 U10041 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n8511), .Z(n8446) );
  NAND2_X1 U10042 ( .A1(n8446), .A2(SI_5_), .ZN(n8449) );
  INV_X1 U10043 ( .A(n8446), .ZN(n8447) );
  INV_X1 U10044 ( .A(SI_5_), .ZN(n10152) );
  NAND2_X1 U10045 ( .A1(n8447), .A2(n10152), .ZN(n8448) );
  MUX2_X1 U10046 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n8511), .Z(n8450) );
  NAND2_X1 U10047 ( .A1(n8450), .A2(SI_6_), .ZN(n8452) );
  OAI21_X1 U10048 ( .B1(n8450), .B2(SI_6_), .A(n8452), .ZN(n8451) );
  INV_X1 U10049 ( .A(n8451), .ZN(n8671) );
  MUX2_X1 U10050 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n8511), .Z(n8453) );
  NAND2_X1 U10051 ( .A1(n8453), .A2(SI_7_), .ZN(n8457) );
  INV_X1 U10052 ( .A(n8453), .ZN(n8454) );
  NAND2_X1 U10053 ( .A1(n8454), .A2(n10148), .ZN(n8455) );
  NAND2_X1 U10054 ( .A1(n8457), .A2(n8455), .ZN(n8688) );
  INV_X1 U10055 ( .A(n8688), .ZN(n8456) );
  MUX2_X1 U10056 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n8511), .Z(n8458) );
  NAND2_X1 U10057 ( .A1(n8458), .A2(SI_8_), .ZN(n8460) );
  OAI21_X1 U10058 ( .B1(n8458), .B2(SI_8_), .A(n8460), .ZN(n8459) );
  INV_X1 U10059 ( .A(n8459), .ZN(n8710) );
  MUX2_X1 U10060 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n8511), .Z(n8461) );
  INV_X1 U10061 ( .A(n8730), .ZN(n8462) );
  MUX2_X1 U10062 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n8511), .Z(n8464) );
  INV_X1 U10063 ( .A(n8464), .ZN(n8465) );
  NAND2_X1 U10064 ( .A1(n8465), .A2(n14440), .ZN(n8466) );
  NAND2_X1 U10065 ( .A1(n8468), .A2(n8466), .ZN(n8749) );
  INV_X1 U10066 ( .A(n8749), .ZN(n8467) );
  MUX2_X1 U10067 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n8511), .Z(n8469) );
  XNOR2_X1 U10068 ( .A(n8469), .B(SI_11_), .ZN(n8769) );
  INV_X1 U10069 ( .A(n8469), .ZN(n8470) );
  MUX2_X1 U10070 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n8511), .Z(n8471) );
  XNOR2_X1 U10071 ( .A(n8471), .B(n14236), .ZN(n8788) );
  INV_X1 U10072 ( .A(n8471), .ZN(n8472) );
  NAND2_X1 U10073 ( .A1(n8472), .A2(n14236), .ZN(n8473) );
  MUX2_X1 U10074 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n8511), .Z(n8475) );
  OAI21_X1 U10075 ( .B1(n8475), .B2(SI_13_), .A(n8476), .ZN(n8811) );
  MUX2_X1 U10076 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n8511), .Z(n8477) );
  XNOR2_X1 U10077 ( .A(n8477), .B(SI_14_), .ZN(n8829) );
  INV_X1 U10078 ( .A(n8477), .ZN(n8478) );
  MUX2_X1 U10079 ( .A(n10650), .B(n10643), .S(n8511), .Z(n8479) );
  NAND2_X1 U10080 ( .A1(n8480), .A2(n14429), .ZN(n8481) );
  MUX2_X1 U10081 ( .A(n11012), .B(n10889), .S(n10468), .Z(n8867) );
  INV_X2 U10082 ( .A(n8511), .ZN(n10165) );
  MUX2_X1 U10083 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n10468), .Z(n8483) );
  MUX2_X1 U10084 ( .A(n11473), .B(n11495), .S(n10468), .Z(n8902) );
  MUX2_X1 U10085 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10468), .Z(n8488) );
  INV_X1 U10086 ( .A(n8488), .ZN(n8489) );
  NAND2_X1 U10087 ( .A1(n8489), .A2(n14424), .ZN(n8490) );
  MUX2_X1 U10088 ( .A(n13177), .B(n12045), .S(n10468), .Z(n8934) );
  XNOR2_X1 U10089 ( .A(n8934), .B(SI_20_), .ZN(n8491) );
  XNOR2_X1 U10090 ( .A(n8936), .B(n8491), .ZN(n13176) );
  NAND2_X1 U10091 ( .A1(n8570), .A2(n8492), .ZN(n8616) );
  INV_X1 U10092 ( .A(n8616), .ZN(n8494) );
  NAND2_X1 U10093 ( .A1(n8494), .A2(n8493), .ZN(n8633) );
  INV_X1 U10094 ( .A(n8633), .ZN(n8504) );
  NOR2_X1 U10095 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8498) );
  NOR2_X2 U10096 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n8496) );
  NOR2_X2 U10097 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n8495) );
  NAND4_X1 U10098 ( .A1(n8498), .A2(n8497), .A3(n8496), .A4(n8495), .ZN(n8798)
         );
  NAND4_X1 U10099 ( .A1(n8501), .A2(n8831), .A3(n8500), .A4(n8499), .ZN(n8502)
         );
  NOR2_X1 U10100 ( .A1(n8798), .A2(n8502), .ZN(n8503) );
  NOR2_X1 U10101 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n8506) );
  NOR2_X1 U10102 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n8505) );
  AND2_X1 U10103 ( .A1(n8506), .A2(n8505), .ZN(n8507) );
  XNOR2_X2 U10104 ( .A(n8510), .B(n8509), .ZN(n15119) );
  NAND2_X2 U10105 ( .A1(n15115), .A2(n15119), .ZN(n8802) );
  INV_X4 U10106 ( .A(n9321), .ZN(n9356) );
  NAND2_X1 U10107 ( .A1(n13176), .A2(n9356), .ZN(n8513) );
  OR2_X1 U10108 ( .A1(n9357), .A2(n12045), .ZN(n8512) );
  NAND2_X1 U10109 ( .A1(n8517), .A2(n8528), .ZN(n9101) );
  NAND2_X1 U10110 ( .A1(n9101), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8518) );
  XNOR2_X1 U10111 ( .A(n8518), .B(P2_IR_REG_22__SCAN_IN), .ZN(n9156) );
  INV_X1 U10112 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8520) );
  NAND2_X1 U10113 ( .A1(n8906), .A2(n8520), .ZN(n8521) );
  AND2_X1 U10114 ( .A1(n8519), .A2(n12727), .ZN(n8530) );
  INV_X1 U10115 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8523) );
  INV_X1 U10116 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8797) );
  AOI21_X1 U10117 ( .B1(n8524), .B2(n8523), .A(n8797), .ZN(n8525) );
  XNOR2_X1 U10118 ( .A(n15053), .B(n9075), .ZN(n8930) );
  NAND2_X1 U10119 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n8659) );
  INV_X1 U10120 ( .A(n8659), .ZN(n8531) );
  NAND2_X1 U10121 ( .A1(n8531), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8678) );
  INV_X1 U10122 ( .A(n8678), .ZN(n8532) );
  NAND2_X1 U10123 ( .A1(n8532), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8697) );
  INV_X1 U10124 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8696) );
  AND2_X1 U10125 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_13__SCAN_IN), 
        .ZN(n8534) );
  INV_X1 U10126 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8857) );
  INV_X1 U10127 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n12534) );
  INV_X1 U10128 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8555) );
  INV_X1 U10129 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n14664) );
  NAND2_X1 U10130 ( .A1(n8557), .A2(n14664), .ZN(n8538) );
  NAND2_X1 U10131 ( .A1(n8943), .A2(n8538), .ZN(n14957) );
  XNOR2_X2 U10132 ( .A(n8540), .B(n15106), .ZN(n12730) );
  NAND2_X2 U10133 ( .A1(n8545), .A2(n8544), .ZN(n8969) );
  INV_X1 U10134 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U10135 ( .A1(n8544), .A2(n15114), .ZN(n8592) );
  INV_X2 U10136 ( .A(n9327), .ZN(n9343) );
  NAND2_X1 U10137 ( .A1(n9343), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U10138 ( .A1(n9342), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8546) );
  OAI211_X1 U10139 ( .C1(n8548), .C2(n9346), .A(n8547), .B(n8546), .ZN(n8549)
         );
  INV_X1 U10140 ( .A(n8549), .ZN(n8550) );
  OAI21_X1 U10141 ( .B1(n14957), .B2(n9341), .A(n8550), .ZN(n14716) );
  NAND2_X1 U10142 ( .A1(n14716), .A2(n14884), .ZN(n8931) );
  XNOR2_X1 U10143 ( .A(n8930), .B(n8931), .ZN(n14662) );
  XNOR2_X1 U10144 ( .A(n8552), .B(n8551), .ZN(n13153) );
  NAND2_X1 U10145 ( .A1(n13153), .A2(n9356), .ZN(n8554) );
  INV_X2 U10146 ( .A(n8802), .ZN(n10271) );
  AOI22_X1 U10147 ( .A1(n8910), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n11851), 
        .B2(n10271), .ZN(n8553) );
  XNOR2_X1 U10148 ( .A(n15057), .B(n9075), .ZN(n8564) );
  NAND2_X1 U10149 ( .A1(n8916), .A2(n8555), .ZN(n8556) );
  NAND2_X1 U10150 ( .A1(n8557), .A2(n8556), .ZN(n14971) );
  OR2_X1 U10151 ( .A1(n14971), .A2(n8969), .ZN(n8563) );
  INV_X1 U10152 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8560) );
  NAND2_X1 U10153 ( .A1(n8894), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8559) );
  NAND2_X1 U10154 ( .A1(n9342), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8558) );
  OAI211_X1 U10155 ( .C1(n9327), .C2(n8560), .A(n8559), .B(n8558), .ZN(n8561)
         );
  INV_X1 U10156 ( .A(n8561), .ZN(n8562) );
  NAND2_X1 U10157 ( .A1(n8563), .A2(n8562), .ZN(n14717) );
  AND2_X1 U10158 ( .A1(n14717), .A2(n14986), .ZN(n8565) );
  NAND2_X1 U10159 ( .A1(n8564), .A2(n8565), .ZN(n8929) );
  INV_X1 U10160 ( .A(n8564), .ZN(n14661) );
  INV_X1 U10161 ( .A(n8565), .ZN(n8566) );
  NAND2_X1 U10162 ( .A1(n14661), .A2(n8566), .ZN(n8567) );
  AND2_X1 U10163 ( .A1(n8929), .A2(n8567), .ZN(n14175) );
  NAND2_X1 U10164 ( .A1(n8614), .A2(SI_2_), .ZN(n8609) );
  NAND2_X1 U10165 ( .A1(n10494), .A2(n9356), .ZN(n8572) );
  INV_X1 U10166 ( .A(n8570), .ZN(n8584) );
  NAND2_X1 U10167 ( .A1(n8584), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8571) );
  XNOR2_X1 U10168 ( .A(n8571), .B(P2_IR_REG_2__SCAN_IN), .ZN(n10282) );
  XNOR2_X1 U10169 ( .A(n10716), .B(n9075), .ZN(n8604) );
  INV_X1 U10170 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10256) );
  OR2_X1 U10171 ( .A1(n9327), .A2(n10256), .ZN(n8577) );
  INV_X1 U10172 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n8573) );
  OR2_X1 U10173 ( .A1(n9346), .A2(n8573), .ZN(n8576) );
  INV_X1 U10174 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10708) );
  OR2_X1 U10175 ( .A1(n8969), .A2(n10708), .ZN(n8574) );
  NAND2_X1 U10176 ( .A1(n14734), .A2(n14884), .ZN(n8605) );
  XNOR2_X1 U10177 ( .A(n8604), .B(n8605), .ZN(n10712) );
  INV_X1 U10178 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10280) );
  INV_X1 U10179 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n8578) );
  OR2_X1 U10180 ( .A1(n8592), .A2(n8578), .ZN(n8581) );
  INV_X1 U10181 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8579) );
  NAND2_X1 U10182 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8583) );
  MUX2_X1 U10183 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8583), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8585) );
  NAND2_X1 U10184 ( .A1(n8585), .A2(n8584), .ZN(n16045) );
  INV_X1 U10185 ( .A(n8586), .ZN(n8587) );
  NAND2_X1 U10186 ( .A1(n8588), .A2(n8587), .ZN(n8589) );
  NAND2_X1 U10187 ( .A1(n8590), .A2(n8589), .ZN(n10467) );
  OR2_X1 U10188 ( .A1(n9321), .A2(n10467), .ZN(n8591) );
  XNOR2_X1 U10189 ( .A(n16420), .B(n8598), .ZN(n10710) );
  XNOR2_X1 U10190 ( .A(n8600), .B(n10710), .ZN(n14208) );
  INV_X1 U10191 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10594) );
  INV_X1 U10192 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10590) );
  INV_X1 U10193 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10589) );
  OR2_X1 U10194 ( .A1(n8592), .A2(n10589), .ZN(n8594) );
  NAND2_X1 U10195 ( .A1(n8894), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8593) );
  INV_X1 U10196 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10591) );
  NAND2_X1 U10197 ( .A1(n8511), .A2(SI_0_), .ZN(n8597) );
  XNOR2_X1 U10198 ( .A(n8597), .B(n9481), .ZN(n15134) );
  MUX2_X1 U10199 ( .A(n10591), .B(n15134), .S(n8802), .Z(n10660) );
  AND2_X1 U10200 ( .A1(n14737), .A2(n8032), .ZN(n14202) );
  AOI21_X1 U10201 ( .B1(n14202), .B2(n14873), .A(n14201), .ZN(n8599) );
  INV_X1 U10202 ( .A(n10710), .ZN(n8601) );
  NAND2_X1 U10203 ( .A1(n8601), .A2(n8600), .ZN(n8602) );
  NAND2_X1 U10204 ( .A1(n10711), .A2(n8602), .ZN(n8603) );
  NAND2_X1 U10205 ( .A1(n10712), .A2(n8603), .ZN(n10718) );
  INV_X1 U10206 ( .A(n8604), .ZN(n8606) );
  NAND2_X1 U10207 ( .A1(n8606), .A2(n8605), .ZN(n8607) );
  NAND2_X1 U10208 ( .A1(n10718), .A2(n8607), .ZN(n14167) );
  AND2_X1 U10209 ( .A1(n8609), .A2(n8608), .ZN(n8610) );
  NAND2_X1 U10210 ( .A1(n8611), .A2(n8610), .ZN(n8615) );
  OAI21_X1 U10211 ( .B1(n8614), .B2(n8613), .A(n8612), .ZN(n8630) );
  AND2_X1 U10212 ( .A1(n8615), .A2(n8630), .ZN(n10516) );
  NAND2_X1 U10213 ( .A1(n10516), .A2(n9356), .ZN(n8619) );
  NAND2_X1 U10214 ( .A1(n8616), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8617) );
  XNOR2_X1 U10215 ( .A(n8617), .B(P2_IR_REG_3__SCAN_IN), .ZN(n14745) );
  AOI22_X1 U10216 ( .A1(n8910), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n10271), 
        .B2(n14745), .ZN(n8618) );
  NAND2_X1 U10217 ( .A1(n8619), .A2(n8618), .ZN(n14170) );
  XNOR2_X1 U10218 ( .A(n14170), .B(n9075), .ZN(n10667) );
  NAND2_X1 U10219 ( .A1(n8894), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8624) );
  INV_X1 U10220 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10285) );
  INV_X1 U10221 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10258) );
  OR2_X1 U10222 ( .A1(n8592), .A2(n10258), .ZN(n8622) );
  OR2_X1 U10223 ( .A1(n8969), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8621) );
  AND2_X1 U10224 ( .A1(n14733), .A2(n14873), .ZN(n8625) );
  NAND2_X1 U10225 ( .A1(n10667), .A2(n8625), .ZN(n8645) );
  INV_X1 U10226 ( .A(n10667), .ZN(n8627) );
  INV_X1 U10227 ( .A(n8625), .ZN(n8626) );
  NAND2_X1 U10228 ( .A1(n8627), .A2(n8626), .ZN(n8628) );
  NAND2_X1 U10229 ( .A1(n8645), .A2(n8628), .ZN(n14166) );
  OR2_X2 U10230 ( .A1(n14167), .A2(n14166), .ZN(n14168) );
  NAND2_X1 U10231 ( .A1(n8630), .A2(n8629), .ZN(n8632) );
  XNOR2_X1 U10232 ( .A(n8631), .B(n8632), .ZN(n10754) );
  NAND2_X1 U10233 ( .A1(n10754), .A2(n9356), .ZN(n8638) );
  NAND2_X1 U10234 ( .A1(n8634), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8635) );
  MUX2_X1 U10235 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8635), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8636) );
  NOR2_X1 U10236 ( .A1(n8634), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8800) );
  INV_X1 U10237 ( .A(n8800), .ZN(n8654) );
  NAND2_X1 U10238 ( .A1(n8636), .A2(n8654), .ZN(n10287) );
  INV_X1 U10239 ( .A(n10287), .ZN(n16071) );
  AOI22_X1 U10240 ( .A1(n8910), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n10271), 
        .B2(n16071), .ZN(n8637) );
  NAND2_X1 U10241 ( .A1(n8638), .A2(n8637), .ZN(n10998) );
  XNOR2_X1 U10242 ( .A(n10998), .B(n9075), .ZN(n8647) );
  NAND2_X1 U10243 ( .A1(n9342), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8644) );
  INV_X1 U10244 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n8639) );
  OR2_X1 U10245 ( .A1(n9327), .A2(n8639), .ZN(n8643) );
  OAI21_X1 U10246 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n8659), .ZN(n16472) );
  OR2_X1 U10247 ( .A1(n8969), .A2(n16472), .ZN(n8642) );
  INV_X1 U10248 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n8640) );
  OR2_X1 U10249 ( .A1(n9346), .A2(n8640), .ZN(n8641) );
  NAND4_X1 U10250 ( .A1(n8644), .A2(n8643), .A3(n8642), .A4(n8641), .ZN(n14732) );
  NAND2_X1 U10251 ( .A1(n14732), .A2(n14884), .ZN(n8648) );
  XNOR2_X1 U10252 ( .A(n8647), .B(n8648), .ZN(n10666) );
  AND2_X1 U10253 ( .A1(n10666), .A2(n8645), .ZN(n8646) );
  INV_X1 U10254 ( .A(n8647), .ZN(n10721) );
  NAND2_X1 U10255 ( .A1(n10721), .A2(n8648), .ZN(n8649) );
  OR2_X1 U10256 ( .A1(n8651), .A2(n8650), .ZN(n8652) );
  NAND2_X1 U10257 ( .A1(n10784), .A2(n9356), .ZN(n8657) );
  NAND2_X1 U10258 ( .A1(n8654), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8653) );
  MUX2_X1 U10259 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8653), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n8655) );
  AND2_X1 U10260 ( .A1(n8655), .A2(n8690), .ZN(n14756) );
  AOI22_X1 U10261 ( .A1(n8910), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n10271), 
        .B2(n14756), .ZN(n8656) );
  XNOR2_X1 U10262 ( .A(n11802), .B(n9075), .ZN(n8667) );
  NAND2_X1 U10263 ( .A1(n9343), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8665) );
  INV_X1 U10264 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10289) );
  OR2_X1 U10265 ( .A1(n8620), .A2(n10289), .ZN(n8664) );
  INV_X1 U10266 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U10267 ( .A1(n8659), .A2(n8658), .ZN(n8660) );
  NAND2_X1 U10268 ( .A1(n8678), .A2(n8660), .ZN(n11799) );
  OR2_X1 U10269 ( .A1(n9341), .A2(n11799), .ZN(n8663) );
  INV_X1 U10270 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n8661) );
  OR2_X1 U10271 ( .A1(n9346), .A2(n8661), .ZN(n8662) );
  NAND4_X1 U10272 ( .A1(n8665), .A2(n8664), .A3(n8663), .A4(n8662), .ZN(n14731) );
  NAND2_X1 U10273 ( .A1(n14731), .A2(n14884), .ZN(n8668) );
  XNOR2_X1 U10274 ( .A(n8667), .B(n8668), .ZN(n10722) );
  INV_X1 U10275 ( .A(n8667), .ZN(n8669) );
  NAND2_X1 U10276 ( .A1(n8669), .A2(n8668), .ZN(n8670) );
  OR2_X1 U10277 ( .A1(n8672), .A2(n8671), .ZN(n8673) );
  NAND2_X1 U10278 ( .A1(n8690), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8675) );
  XNOR2_X1 U10279 ( .A(n8675), .B(P2_IR_REG_6__SCAN_IN), .ZN(n14769) );
  AOI22_X1 U10280 ( .A1(n8910), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n10271), 
        .B2(n14769), .ZN(n8676) );
  XNOR2_X1 U10281 ( .A(n11934), .B(n9075), .ZN(n10848) );
  NAND2_X1 U10282 ( .A1(n8894), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8683) );
  INV_X1 U10283 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10292) );
  OR2_X1 U10284 ( .A1(n8620), .A2(n10292), .ZN(n8682) );
  INV_X1 U10285 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8677) );
  NAND2_X1 U10286 ( .A1(n8678), .A2(n8677), .ZN(n8679) );
  NAND2_X1 U10287 ( .A1(n8697), .A2(n8679), .ZN(n11930) );
  OR2_X1 U10288 ( .A1(n8969), .A2(n11930), .ZN(n8681) );
  INV_X1 U10289 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11931) );
  OR2_X1 U10290 ( .A1(n9327), .A2(n11931), .ZN(n8680) );
  NAND4_X1 U10291 ( .A1(n8683), .A2(n8682), .A3(n8681), .A4(n8680), .ZN(n14730) );
  AND2_X1 U10292 ( .A1(n14730), .A2(n14986), .ZN(n8684) );
  NAND2_X1 U10293 ( .A1(n10848), .A2(n8684), .ZN(n8704) );
  INV_X1 U10294 ( .A(n10848), .ZN(n8686) );
  INV_X1 U10295 ( .A(n8684), .ZN(n8685) );
  NAND2_X1 U10296 ( .A1(n8686), .A2(n8685), .ZN(n8687) );
  NAND2_X1 U10297 ( .A1(n8704), .A2(n8687), .ZN(n11047) );
  NAND2_X1 U10298 ( .A1(n11060), .A2(n9356), .ZN(n8695) );
  INV_X1 U10299 ( .A(n8690), .ZN(n8692) );
  INV_X1 U10300 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U10301 ( .A1(n8692), .A2(n8691), .ZN(n8714) );
  NAND2_X1 U10302 ( .A1(n8714), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8693) );
  XNOR2_X1 U10303 ( .A(n8693), .B(P2_IR_REG_7__SCAN_IN), .ZN(n14783) );
  AOI22_X1 U10304 ( .A1(n8910), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n10271), 
        .B2(n14783), .ZN(n8694) );
  XNOR2_X1 U10305 ( .A(n11548), .B(n9075), .ZN(n8706) );
  NAND2_X1 U10306 ( .A1(n9342), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8703) );
  INV_X1 U10307 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10264) );
  OR2_X1 U10308 ( .A1(n9327), .A2(n10264), .ZN(n8702) );
  NAND2_X1 U10309 ( .A1(n8697), .A2(n8696), .ZN(n8698) );
  NAND2_X1 U10310 ( .A1(n8719), .A2(n8698), .ZN(n16510) );
  OR2_X1 U10311 ( .A1(n9341), .A2(n16510), .ZN(n8701) );
  INV_X1 U10312 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8699) );
  OR2_X1 U10313 ( .A1(n9346), .A2(n8699), .ZN(n8700) );
  NAND4_X1 U10314 ( .A1(n8703), .A2(n8702), .A3(n8701), .A4(n8700), .ZN(n14729) );
  NAND2_X1 U10315 ( .A1(n14729), .A2(n14884), .ZN(n8707) );
  XNOR2_X1 U10316 ( .A(n8706), .B(n8707), .ZN(n10850) );
  AND2_X1 U10317 ( .A1(n10850), .A2(n8704), .ZN(n8705) );
  INV_X1 U10318 ( .A(n8706), .ZN(n8708) );
  NAND2_X1 U10319 ( .A1(n8708), .A2(n8707), .ZN(n8709) );
  NAND2_X1 U10320 ( .A1(n10855), .A2(n8709), .ZN(n11157) );
  OR2_X1 U10321 ( .A1(n8711), .A2(n8710), .ZN(n8712) );
  NAND2_X1 U10322 ( .A1(n8713), .A2(n8712), .ZN(n11290) );
  OR2_X1 U10323 ( .A1(n11290), .A2(n9321), .ZN(n8717) );
  NAND2_X1 U10324 ( .A1(n8732), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8715) );
  XNOR2_X1 U10325 ( .A(n8715), .B(P2_IR_REG_8__SCAN_IN), .ZN(n14797) );
  AOI22_X1 U10326 ( .A1(n8910), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n10271), 
        .B2(n14797), .ZN(n8716) );
  XNOR2_X1 U10327 ( .A(n12034), .B(n14190), .ZN(n8726) );
  NAND2_X1 U10328 ( .A1(n9343), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8725) );
  INV_X1 U10329 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10298) );
  OR2_X1 U10330 ( .A1(n8620), .A2(n10298), .ZN(n8724) );
  NAND2_X1 U10331 ( .A1(n8719), .A2(n8718), .ZN(n8720) );
  NAND2_X1 U10332 ( .A1(n8736), .A2(n8720), .ZN(n12038) );
  OR2_X1 U10333 ( .A1(n9341), .A2(n12038), .ZN(n8723) );
  INV_X1 U10334 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n8721) );
  OR2_X1 U10335 ( .A1(n9346), .A2(n8721), .ZN(n8722) );
  NAND4_X1 U10336 ( .A1(n8725), .A2(n8724), .A3(n8723), .A4(n8722), .ZN(n14728) );
  NAND2_X1 U10337 ( .A1(n14728), .A2(n14884), .ZN(n8727) );
  AND2_X1 U10338 ( .A1(n8726), .A2(n8727), .ZN(n11153) );
  INV_X1 U10339 ( .A(n8726), .ZN(n8729) );
  INV_X1 U10340 ( .A(n8727), .ZN(n8728) );
  NAND2_X1 U10341 ( .A1(n8729), .A2(n8728), .ZN(n11154) );
  XNOR2_X1 U10342 ( .A(n8731), .B(n8730), .ZN(n11416) );
  NAND2_X1 U10343 ( .A1(n11416), .A2(n9356), .ZN(n8734) );
  NAND2_X1 U10344 ( .A1(n8790), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8751) );
  XNOR2_X1 U10345 ( .A(n8751), .B(P2_IR_REG_9__SCAN_IN), .ZN(n16151) );
  AOI22_X1 U10346 ( .A1(n10271), .A2(n16151), .B1(n8910), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n8733) );
  XNOR2_X1 U10347 ( .A(n12095), .B(n14190), .ZN(n8743) );
  NAND2_X1 U10348 ( .A1(n9342), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8742) );
  INV_X1 U10349 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n12098) );
  OR2_X1 U10350 ( .A1(n9327), .A2(n12098), .ZN(n8741) );
  NAND2_X1 U10351 ( .A1(n8736), .A2(n8735), .ZN(n8737) );
  NAND2_X1 U10352 ( .A1(n8756), .A2(n8737), .ZN(n12097) );
  OR2_X1 U10353 ( .A1(n9341), .A2(n12097), .ZN(n8740) );
  INV_X1 U10354 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8738) );
  OR2_X1 U10355 ( .A1(n9346), .A2(n8738), .ZN(n8739) );
  NAND4_X1 U10356 ( .A1(n8742), .A2(n8741), .A3(n8740), .A4(n8739), .ZN(n14727) );
  NAND2_X1 U10357 ( .A1(n14727), .A2(n14873), .ZN(n8744) );
  NAND2_X1 U10358 ( .A1(n8743), .A2(n8744), .ZN(n8748) );
  INV_X1 U10359 ( .A(n8743), .ZN(n8746) );
  INV_X1 U10360 ( .A(n8744), .ZN(n8745) );
  NAND2_X1 U10361 ( .A1(n8746), .A2(n8745), .ZN(n8747) );
  NAND2_X1 U10362 ( .A1(n8748), .A2(n8747), .ZN(n11378) );
  OR2_X2 U10363 ( .A1(n11377), .A2(n11378), .ZN(n11375) );
  XNOR2_X1 U10364 ( .A(n8750), .B(n8749), .ZN(n11585) );
  NAND2_X1 U10365 ( .A1(n11585), .A2(n9356), .ZN(n8754) );
  INV_X1 U10366 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8793) );
  NAND2_X1 U10367 ( .A1(n8751), .A2(n8793), .ZN(n8752) );
  NAND2_X1 U10368 ( .A1(n8752), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8771) );
  XNOR2_X1 U10369 ( .A(n8771), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10372) );
  AOI22_X1 U10370 ( .A1(n10372), .A2(n10271), .B1(n8910), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n8753) );
  XNOR2_X1 U10371 ( .A(n12151), .B(n14190), .ZN(n8763) );
  NAND2_X1 U10372 ( .A1(n9342), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8762) );
  INV_X1 U10373 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n12149) );
  OR2_X1 U10374 ( .A1(n9327), .A2(n12149), .ZN(n8761) );
  INV_X1 U10375 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U10376 ( .A1(n8756), .A2(n8755), .ZN(n8757) );
  NAND2_X1 U10377 ( .A1(n8777), .A2(n8757), .ZN(n12148) );
  OR2_X1 U10378 ( .A1(n9341), .A2(n12148), .ZN(n8760) );
  INV_X1 U10379 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n8758) );
  OR2_X1 U10380 ( .A1(n9346), .A2(n8758), .ZN(n8759) );
  NAND4_X1 U10381 ( .A1(n8762), .A2(n8761), .A3(n8760), .A4(n8759), .ZN(n14726) );
  NAND2_X1 U10382 ( .A1(n14726), .A2(n14884), .ZN(n8764) );
  NAND2_X1 U10383 ( .A1(n8763), .A2(n8764), .ZN(n8768) );
  INV_X1 U10384 ( .A(n8763), .ZN(n8766) );
  INV_X1 U10385 ( .A(n8764), .ZN(n8765) );
  NAND2_X1 U10386 ( .A1(n8766), .A2(n8765), .ZN(n8767) );
  AND2_X1 U10387 ( .A1(n8768), .A2(n8767), .ZN(n11461) );
  XNOR2_X1 U10388 ( .A(n8770), .B(n8769), .ZN(n11862) );
  NAND2_X1 U10389 ( .A1(n11862), .A2(n9356), .ZN(n8775) );
  INV_X1 U10390 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n8792) );
  NAND2_X1 U10391 ( .A1(n8771), .A2(n8792), .ZN(n8772) );
  NAND2_X1 U10392 ( .A1(n8772), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8773) );
  XNOR2_X1 U10393 ( .A(n8773), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10576) );
  AOI22_X1 U10394 ( .A1(n10576), .A2(n10271), .B1(n8910), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8774) );
  XNOR2_X1 U10395 ( .A(n12223), .B(n14190), .ZN(n8784) );
  NAND2_X1 U10396 ( .A1(n9342), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8783) );
  INV_X1 U10397 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8776) );
  OR2_X1 U10398 ( .A1(n9327), .A2(n8776), .ZN(n8782) );
  NAND2_X1 U10399 ( .A1(n8777), .A2(n10368), .ZN(n8778) );
  NAND2_X1 U10400 ( .A1(n8820), .A2(n8778), .ZN(n11695) );
  OR2_X1 U10401 ( .A1(n9341), .A2(n11695), .ZN(n8781) );
  INV_X1 U10402 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8779) );
  OR2_X1 U10403 ( .A1(n9346), .A2(n8779), .ZN(n8780) );
  NAND4_X1 U10404 ( .A1(n8783), .A2(n8782), .A3(n8781), .A4(n8780), .ZN(n14725) );
  NAND2_X1 U10405 ( .A1(n14725), .A2(n14873), .ZN(n8785) );
  XNOR2_X1 U10406 ( .A(n8784), .B(n8785), .ZN(n11694) );
  INV_X1 U10407 ( .A(n8784), .ZN(n8787) );
  INV_X1 U10408 ( .A(n8785), .ZN(n8786) );
  XNOR2_X1 U10409 ( .A(n8789), .B(n8788), .ZN(n11959) );
  NAND2_X1 U10410 ( .A1(n11959), .A2(n9356), .ZN(n8805) );
  INV_X1 U10411 ( .A(n8790), .ZN(n8795) );
  INV_X1 U10412 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n8791) );
  AND3_X1 U10413 ( .A1(n8793), .A2(n8792), .A3(n8791), .ZN(n8794) );
  AOI21_X1 U10414 ( .B1(n8795), .B2(n8794), .A(n8797), .ZN(n8796) );
  MUX2_X1 U10415 ( .A(n8797), .B(n8796), .S(P2_IR_REG_12__SCAN_IN), .Z(n8801)
         );
  INV_X1 U10416 ( .A(n8798), .ZN(n8799) );
  AND2_X1 U10417 ( .A1(n8800), .A2(n8799), .ZN(n8832) );
  OAI22_X1 U10418 ( .A1(n16126), .A2(n8802), .B1(n9357), .B2(n10248), .ZN(
        n8803) );
  INV_X1 U10419 ( .A(n8803), .ZN(n8804) );
  XNOR2_X1 U10420 ( .A(n16606), .B(n9075), .ZN(n14626) );
  NAND2_X1 U10421 ( .A1(n9343), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8810) );
  INV_X1 U10422 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10569) );
  OR2_X1 U10423 ( .A1(n8620), .A2(n10569), .ZN(n8809) );
  INV_X1 U10424 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8819) );
  XNOR2_X1 U10425 ( .A(n8820), .B(n8819), .ZN(n14631) );
  OR2_X1 U10426 ( .A1(n9341), .A2(n14631), .ZN(n8808) );
  INV_X1 U10427 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8806) );
  OR2_X1 U10428 ( .A1(n9346), .A2(n8806), .ZN(n8807) );
  NAND4_X1 U10429 ( .A1(n8810), .A2(n8809), .A3(n8808), .A4(n8807), .ZN(n14724) );
  AND2_X1 U10430 ( .A1(n14724), .A2(n14986), .ZN(n14627) );
  AND2_X1 U10431 ( .A1(n14626), .A2(n14627), .ZN(n14624) );
  XNOR2_X1 U10432 ( .A(n8812), .B(n8279), .ZN(n11999) );
  NAND2_X1 U10433 ( .A1(n11999), .A2(n9356), .ZN(n8816) );
  INV_X1 U10434 ( .A(n8832), .ZN(n8813) );
  NAND2_X1 U10435 ( .A1(n8813), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8814) );
  XNOR2_X1 U10436 ( .A(n8814), .B(P2_IR_REG_13__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U10437 ( .A1(n8910), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n10271), 
        .B2(n10572), .ZN(n8815) );
  XNOR2_X1 U10438 ( .A(n12427), .B(n14190), .ZN(n12133) );
  NAND2_X1 U10439 ( .A1(n9342), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8825) );
  INV_X1 U10440 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8817) );
  OR2_X1 U10441 ( .A1(n9346), .A2(n8817), .ZN(n8824) );
  INV_X1 U10442 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8818) );
  OAI21_X1 U10443 ( .B1(n8820), .B2(n8819), .A(n8818), .ZN(n8821) );
  NAND2_X1 U10444 ( .A1(n8837), .A2(n8821), .ZN(n12274) );
  OR2_X1 U10445 ( .A1(n9341), .A2(n12274), .ZN(n8823) );
  INV_X1 U10446 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10691) );
  OR2_X1 U10447 ( .A1(n9327), .A2(n10691), .ZN(n8822) );
  NAND4_X1 U10448 ( .A1(n8825), .A2(n8824), .A3(n8823), .A4(n8822), .ZN(n14723) );
  NAND2_X1 U10449 ( .A1(n14723), .A2(n14873), .ZN(n8827) );
  XNOR2_X1 U10450 ( .A(n12133), .B(n8827), .ZN(n12088) );
  AOI21_X1 U10451 ( .B1(n14629), .B2(n14627), .A(n12088), .ZN(n8826) );
  NAND2_X1 U10452 ( .A1(n12133), .A2(n8827), .ZN(n8828) );
  XNOR2_X1 U10453 ( .A(n8830), .B(n8829), .ZN(n12312) );
  NAND2_X1 U10454 ( .A1(n12312), .A2(n9356), .ZN(n8835) );
  NAND2_X1 U10455 ( .A1(n8832), .A2(n8831), .ZN(n8851) );
  NAND2_X1 U10456 ( .A1(n8851), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8833) );
  XNOR2_X1 U10457 ( .A(n8833), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U10458 ( .A1(n8910), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n10271), 
        .B2(n11837), .ZN(n8834) );
  XNOR2_X1 U10459 ( .A(n12566), .B(n9075), .ZN(n8845) );
  NAND2_X1 U10460 ( .A1(n8837), .A2(n12129), .ZN(n8838) );
  AND2_X1 U10461 ( .A1(n8858), .A2(n8838), .ZN(n12378) );
  NAND2_X1 U10462 ( .A1(n8836), .A2(n12378), .ZN(n8844) );
  INV_X1 U10463 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8839) );
  OR2_X1 U10464 ( .A1(n8620), .A2(n8839), .ZN(n8843) );
  INV_X1 U10465 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8840) );
  OR2_X1 U10466 ( .A1(n9346), .A2(n8840), .ZN(n8842) );
  INV_X1 U10467 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11840) );
  OR2_X1 U10468 ( .A1(n9327), .A2(n11840), .ZN(n8841) );
  NAND4_X1 U10469 ( .A1(n8844), .A2(n8843), .A3(n8842), .A4(n8841), .ZN(n14722) );
  NAND2_X1 U10470 ( .A1(n14722), .A2(n14873), .ZN(n8846) );
  XNOR2_X1 U10471 ( .A(n8845), .B(n8846), .ZN(n12132) );
  INV_X1 U10472 ( .A(n8845), .ZN(n8847) );
  NAND2_X1 U10473 ( .A1(n8847), .A2(n8846), .ZN(n8848) );
  XNOR2_X1 U10474 ( .A(n8850), .B(n8849), .ZN(n12402) );
  NAND2_X1 U10475 ( .A1(n12402), .A2(n9356), .ZN(n8854) );
  OAI21_X1 U10476 ( .B1(n8851), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8852) );
  XNOR2_X1 U10477 ( .A(n8852), .B(P2_IR_REG_15__SCAN_IN), .ZN(n16079) );
  AOI22_X1 U10478 ( .A1(n8910), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n10271), 
        .B2(n16079), .ZN(n8853) );
  XNOR2_X1 U10479 ( .A(n15078), .B(n9075), .ZN(n8863) );
  INV_X1 U10480 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8856) );
  NAND2_X1 U10481 ( .A1(n9342), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8855) );
  OAI21_X1 U10482 ( .B1(n8856), .B2(n9327), .A(n8855), .ZN(n8862) );
  NAND2_X1 U10483 ( .A1(n8858), .A2(n8857), .ZN(n8859) );
  NAND2_X1 U10484 ( .A1(n8877), .A2(n8859), .ZN(n12606) );
  NAND2_X1 U10485 ( .A1(n8894), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8860) );
  OAI21_X1 U10486 ( .B1(n12606), .B2(n9341), .A(n8860), .ZN(n8861) );
  AND2_X1 U10487 ( .A1(n14721), .A2(n14986), .ZN(n8864) );
  NAND2_X1 U10488 ( .A1(n8863), .A2(n8864), .ZN(n8882) );
  INV_X1 U10489 ( .A(n8863), .ZN(n12627) );
  INV_X1 U10490 ( .A(n8864), .ZN(n8865) );
  NAND2_X1 U10491 ( .A1(n12627), .A2(n8865), .ZN(n8866) );
  NAND2_X1 U10492 ( .A1(n8882), .A2(n8866), .ZN(n12608) );
  OR2_X2 U10493 ( .A1(n12609), .A2(n12608), .ZN(n12607) );
  NAND2_X1 U10494 ( .A1(n8868), .A2(n8867), .ZN(n8869) );
  NAND2_X1 U10495 ( .A1(n13109), .A2(n9356), .ZN(n8875) );
  INV_X1 U10496 ( .A(n8871), .ZN(n8872) );
  NAND2_X1 U10497 ( .A1(n8872), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8873) );
  XNOR2_X1 U10498 ( .A(n8873), .B(P2_IR_REG_16__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U10499 ( .A1(n8910), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n10271), 
        .B2(n11836), .ZN(n8874) );
  XNOR2_X1 U10500 ( .A(n15073), .B(n9075), .ZN(n8884) );
  INV_X1 U10501 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8881) );
  INV_X1 U10502 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8876) );
  NAND2_X1 U10503 ( .A1(n8877), .A2(n8876), .ZN(n8878) );
  NAND2_X1 U10504 ( .A1(n8892), .A2(n8878), .ZN(n12633) );
  OR2_X1 U10505 ( .A1(n12633), .A2(n9341), .ZN(n8880) );
  AOI22_X1 U10506 ( .A1(n9343), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n9342), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n8879) );
  OAI211_X1 U10507 ( .C1(n9346), .C2(n8881), .A(n8880), .B(n8879), .ZN(n14720)
         );
  NAND2_X1 U10508 ( .A1(n14720), .A2(n14873), .ZN(n8885) );
  XNOR2_X1 U10509 ( .A(n8884), .B(n8885), .ZN(n12638) );
  AND2_X1 U10510 ( .A1(n12638), .A2(n8882), .ZN(n8883) );
  NAND2_X2 U10511 ( .A1(n12607), .A2(n8883), .ZN(n12634) );
  INV_X1 U10512 ( .A(n8884), .ZN(n12538) );
  NAND2_X1 U10513 ( .A1(n12538), .A2(n8885), .ZN(n8886) );
  XNOR2_X1 U10514 ( .A(n8888), .B(n8887), .ZN(n13127) );
  NAND2_X1 U10515 ( .A1(n13127), .A2(n9356), .ZN(n8891) );
  NAND2_X1 U10516 ( .A1(n8889), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8907) );
  XNOR2_X1 U10517 ( .A(n8907), .B(P2_IR_REG_17__SCAN_IN), .ZN(n16102) );
  AOI22_X1 U10518 ( .A1(n8910), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n10271), 
        .B2(n16102), .ZN(n8890) );
  XNOR2_X1 U10519 ( .A(n15068), .B(n9075), .ZN(n8898) );
  NAND2_X1 U10520 ( .A1(n8892), .A2(n12534), .ZN(n8893) );
  NAND2_X1 U10521 ( .A1(n8914), .A2(n8893), .ZN(n12654) );
  AOI22_X1 U10522 ( .A1(n9343), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9342), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n8896) );
  NAND2_X1 U10523 ( .A1(n8894), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8895) );
  OAI211_X1 U10524 ( .C1(n12654), .C2(n9341), .A(n8896), .B(n8895), .ZN(n14719) );
  NAND2_X1 U10525 ( .A1(n14719), .A2(n14873), .ZN(n8899) );
  XNOR2_X1 U10526 ( .A(n8898), .B(n8899), .ZN(n12537) );
  INV_X1 U10527 ( .A(n8898), .ZN(n8900) );
  NAND2_X1 U10528 ( .A1(n8900), .A2(n8899), .ZN(n8901) );
  NAND2_X1 U10529 ( .A1(n8903), .A2(n8902), .ZN(n8904) );
  AND2_X1 U10530 ( .A1(n8905), .A2(n8904), .ZN(n13135) );
  NAND2_X1 U10531 ( .A1(n13135), .A2(n9356), .ZN(n8912) );
  NAND2_X1 U10532 ( .A1(n8907), .A2(n8906), .ZN(n8908) );
  NAND2_X1 U10533 ( .A1(n8908), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8909) );
  XNOR2_X1 U10534 ( .A(n8909), .B(P2_IR_REG_18__SCAN_IN), .ZN(n16115) );
  AOI22_X1 U10535 ( .A1(n8910), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n10271), 
        .B2(n16115), .ZN(n8911) );
  XNOR2_X1 U10536 ( .A(n15062), .B(n9075), .ZN(n8923) );
  INV_X1 U10537 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8913) );
  NAND2_X1 U10538 ( .A1(n8914), .A2(n8913), .ZN(n8915) );
  NAND2_X1 U10539 ( .A1(n8916), .A2(n8915), .ZN(n14990) );
  OR2_X1 U10540 ( .A1(n14990), .A2(n8969), .ZN(n8922) );
  INV_X1 U10541 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8919) );
  NAND2_X1 U10542 ( .A1(n9342), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8918) );
  NAND2_X1 U10543 ( .A1(n9343), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8917) );
  OAI211_X1 U10544 ( .C1(n9346), .C2(n8919), .A(n8918), .B(n8917), .ZN(n8920)
         );
  INV_X1 U10545 ( .A(n8920), .ZN(n8921) );
  NAND2_X1 U10546 ( .A1(n8922), .A2(n8921), .ZN(n14718) );
  AND2_X1 U10547 ( .A1(n14718), .A2(n14986), .ZN(n8924) );
  NAND2_X1 U10548 ( .A1(n8923), .A2(n8924), .ZN(n8927) );
  INV_X1 U10549 ( .A(n8923), .ZN(n14178) );
  INV_X1 U10550 ( .A(n8924), .ZN(n8925) );
  NAND2_X1 U10551 ( .A1(n14178), .A2(n8925), .ZN(n8926) );
  NAND2_X1 U10552 ( .A1(n8927), .A2(n8926), .ZN(n14687) );
  NAND2_X1 U10553 ( .A1(n14175), .A2(n8928), .ZN(n14660) );
  INV_X1 U10554 ( .A(n8930), .ZN(n8932) );
  NAND2_X1 U10555 ( .A1(n8932), .A2(n8931), .ZN(n8933) );
  NOR2_X1 U10556 ( .A1(n8937), .A2(SI_20_), .ZN(n8935) );
  NAND2_X1 U10557 ( .A1(n8937), .A2(SI_20_), .ZN(n8938) );
  MUX2_X1 U10558 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10468), .Z(n8959) );
  XNOR2_X1 U10559 ( .A(n8959), .B(SI_21_), .ZN(n8956) );
  XNOR2_X1 U10560 ( .A(n8958), .B(n8956), .ZN(n13182) );
  NAND2_X1 U10561 ( .A1(n13182), .A2(n9356), .ZN(n8940) );
  INV_X1 U10562 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12141) );
  OR2_X1 U10563 ( .A1(n9357), .A2(n12141), .ZN(n8939) );
  XNOR2_X1 U10564 ( .A(n15048), .B(n14190), .ZN(n8951) );
  INV_X1 U10565 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8942) );
  NAND2_X1 U10566 ( .A1(n8943), .A2(n8942), .ZN(n8944) );
  AND2_X1 U10567 ( .A1(n8967), .A2(n8944), .ZN(n14934) );
  NAND2_X1 U10568 ( .A1(n14934), .A2(n8836), .ZN(n8950) );
  INV_X1 U10569 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8947) );
  NAND2_X1 U10570 ( .A1(n9343), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8946) );
  NAND2_X1 U10571 ( .A1(n9342), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8945) );
  OAI211_X1 U10572 ( .C1(n8947), .C2(n9346), .A(n8946), .B(n8945), .ZN(n8948)
         );
  INV_X1 U10573 ( .A(n8948), .ZN(n8949) );
  NAND2_X1 U10574 ( .A1(n8950), .A2(n8949), .ZN(n14912) );
  NAND2_X1 U10575 ( .A1(n14912), .A2(n14873), .ZN(n8952) );
  XNOR2_X1 U10576 ( .A(n8951), .B(n8952), .ZN(n14616) );
  INV_X1 U10577 ( .A(n8951), .ZN(n8954) );
  INV_X1 U10578 ( .A(n8952), .ZN(n8953) );
  NAND2_X1 U10579 ( .A1(n8954), .A2(n8953), .ZN(n8955) );
  INV_X1 U10580 ( .A(SI_22_), .ZN(n14417) );
  MUX2_X1 U10581 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n10468), .Z(n8960) );
  INV_X1 U10582 ( .A(n13203), .ZN(n8961) );
  NAND2_X1 U10583 ( .A1(n8961), .A2(n8256), .ZN(n8962) );
  NAND2_X1 U10584 ( .A1(n8983), .A2(n8962), .ZN(n12299) );
  INV_X1 U10585 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12298) );
  OR2_X1 U10586 ( .A1(n9357), .A2(n12298), .ZN(n8963) );
  XNOR2_X1 U10587 ( .A(n15039), .B(n14190), .ZN(n8977) );
  INV_X1 U10588 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8966) );
  NAND2_X1 U10589 ( .A1(n8967), .A2(n8966), .ZN(n8968) );
  NAND2_X1 U10590 ( .A1(n9004), .A2(n8968), .ZN(n14921) );
  OR2_X1 U10591 ( .A1(n14921), .A2(n8969), .ZN(n8975) );
  INV_X1 U10592 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8972) );
  NAND2_X1 U10593 ( .A1(n9343), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8971) );
  NAND2_X1 U10594 ( .A1(n9342), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8970) );
  OAI211_X1 U10595 ( .C1(n8972), .C2(n9346), .A(n8971), .B(n8970), .ZN(n8973)
         );
  INV_X1 U10596 ( .A(n8973), .ZN(n8974) );
  NAND2_X1 U10597 ( .A1(n8975), .A2(n8974), .ZN(n14715) );
  AND2_X1 U10598 ( .A1(n14715), .A2(n14986), .ZN(n8976) );
  NAND2_X1 U10599 ( .A1(n14672), .A2(n8976), .ZN(n14673) );
  INV_X1 U10600 ( .A(n8977), .ZN(n8978) );
  NAND2_X1 U10601 ( .A1(n8979), .A2(n8978), .ZN(n8980) );
  NAND2_X1 U10602 ( .A1(n14673), .A2(n8980), .ZN(n8994) );
  NAND2_X1 U10603 ( .A1(n8981), .A2(SI_22_), .ZN(n8982) );
  MUX2_X1 U10604 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10468), .Z(n8998) );
  XNOR2_X1 U10605 ( .A(n8998), .B(SI_23_), .ZN(n8996) );
  XNOR2_X1 U10606 ( .A(n8997), .B(n8996), .ZN(n13218) );
  NAND2_X1 U10607 ( .A1(n13218), .A2(n9356), .ZN(n8985) );
  INV_X1 U10608 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n12473) );
  OR2_X1 U10609 ( .A1(n9357), .A2(n12473), .ZN(n8984) );
  XNOR2_X1 U10610 ( .A(n15035), .B(n14190), .ZN(n8992) );
  XNOR2_X1 U10611 ( .A(n8994), .B(n8992), .ZN(n14158) );
  XNOR2_X1 U10612 ( .A(n9004), .B(P2_REG3_REG_23__SCAN_IN), .ZN(n14904) );
  NAND2_X1 U10613 ( .A1(n14904), .A2(n8836), .ZN(n8991) );
  INV_X1 U10614 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8988) );
  NAND2_X1 U10615 ( .A1(n9343), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8987) );
  NAND2_X1 U10616 ( .A1(n9342), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8986) );
  OAI211_X1 U10617 ( .C1(n8988), .C2(n9346), .A(n8987), .B(n8986), .ZN(n8989)
         );
  INV_X1 U10618 ( .A(n8989), .ZN(n8990) );
  NAND2_X1 U10619 ( .A1(n14914), .A2(n14884), .ZN(n14157) );
  INV_X1 U10620 ( .A(n8992), .ZN(n8993) );
  OR2_X1 U10621 ( .A1(n8994), .A2(n8993), .ZN(n8995) );
  NAND2_X1 U10622 ( .A1(n8998), .A2(SI_23_), .ZN(n8999) );
  INV_X1 U10623 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n15993) );
  INV_X1 U10624 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n15132) );
  MUX2_X1 U10625 ( .A(n15993), .B(n15132), .S(n10468), .Z(n9021) );
  XNOR2_X1 U10626 ( .A(n9021), .B(SI_24_), .ZN(n9019) );
  INV_X1 U10627 ( .A(n9019), .ZN(n9000) );
  XNOR2_X1 U10628 ( .A(n9020), .B(n9000), .ZN(n15129) );
  NAND2_X1 U10629 ( .A1(n15129), .A2(n9356), .ZN(n9002) );
  OR2_X1 U10630 ( .A1(n9357), .A2(n15132), .ZN(n9001) );
  XNOR2_X1 U10631 ( .A(n14889), .B(n14190), .ZN(n9014) );
  INV_X1 U10632 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n14161) );
  INV_X1 U10633 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9003) );
  OAI21_X1 U10634 ( .B1(n9004), .B2(n14161), .A(n9003), .ZN(n9007) );
  INV_X1 U10635 ( .A(n9004), .ZN(n9006) );
  AND2_X1 U10636 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .ZN(n9005) );
  INV_X1 U10637 ( .A(n9030), .ZN(n9032) );
  NAND2_X1 U10638 ( .A1(n14887), .A2(n8836), .ZN(n9013) );
  INV_X1 U10639 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9010) );
  NAND2_X1 U10640 ( .A1(n9343), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9009) );
  NAND2_X1 U10641 ( .A1(n9342), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9008) );
  OAI211_X1 U10642 ( .C1(n9010), .C2(n9346), .A(n9009), .B(n9008), .ZN(n9011)
         );
  INV_X1 U10643 ( .A(n9011), .ZN(n9012) );
  NOR2_X1 U10644 ( .A1(n14870), .A2(n14930), .ZN(n9015) );
  NAND2_X1 U10645 ( .A1(n9014), .A2(n9015), .ZN(n9018) );
  INV_X1 U10646 ( .A(n9014), .ZN(n14640) );
  INV_X1 U10647 ( .A(n9015), .ZN(n9016) );
  NAND2_X1 U10648 ( .A1(n14640), .A2(n9016), .ZN(n9017) );
  NAND2_X1 U10649 ( .A1(n9018), .A2(n9017), .ZN(n14654) );
  NAND2_X1 U10650 ( .A1(n9020), .A2(n9019), .ZN(n9024) );
  INV_X1 U10651 ( .A(n9021), .ZN(n9022) );
  NAND2_X1 U10652 ( .A1(n9022), .A2(SI_24_), .ZN(n9023) );
  INV_X1 U10653 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15988) );
  INV_X1 U10654 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n15128) );
  MUX2_X1 U10655 ( .A(n15988), .B(n15128), .S(n8511), .Z(n9025) );
  INV_X1 U10656 ( .A(SI_25_), .ZN(n12349) );
  NAND2_X1 U10657 ( .A1(n9025), .A2(n12349), .ZN(n9047) );
  INV_X1 U10658 ( .A(n9025), .ZN(n9026) );
  NAND2_X1 U10659 ( .A1(n9026), .A2(SI_25_), .ZN(n9027) );
  NAND2_X1 U10660 ( .A1(n9047), .A2(n9027), .ZN(n9045) );
  XNOR2_X1 U10661 ( .A(n9046), .B(n9045), .ZN(n15126) );
  NAND2_X1 U10662 ( .A1(n15126), .A2(n9356), .ZN(n9029) );
  OR2_X1 U10663 ( .A1(n9357), .A2(n15128), .ZN(n9028) );
  XNOR2_X1 U10664 ( .A(n14877), .B(n14190), .ZN(n9040) );
  INV_X1 U10665 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9031) );
  NAND2_X1 U10666 ( .A1(n9032), .A2(n9031), .ZN(n9033) );
  NAND2_X1 U10667 ( .A1(n9054), .A2(n9033), .ZN(n14643) );
  INV_X1 U10668 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9036) );
  NAND2_X1 U10669 ( .A1(n9343), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9035) );
  NAND2_X1 U10670 ( .A1(n9342), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n9034) );
  OAI211_X1 U10671 ( .C1(n9036), .C2(n9346), .A(n9035), .B(n9034), .ZN(n9037)
         );
  INV_X1 U10672 ( .A(n9037), .ZN(n9038) );
  NOR2_X1 U10673 ( .A1(n14695), .A2(n14930), .ZN(n9041) );
  NAND2_X1 U10674 ( .A1(n9040), .A2(n9041), .ZN(n9062) );
  INV_X1 U10675 ( .A(n9040), .ZN(n14696) );
  INV_X1 U10676 ( .A(n9041), .ZN(n9042) );
  NAND2_X1 U10677 ( .A1(n14696), .A2(n9042), .ZN(n9043) );
  AND2_X1 U10678 ( .A1(n9062), .A2(n9043), .ZN(n14638) );
  MUX2_X1 U10679 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n10468), .Z(n9068) );
  XNOR2_X1 U10680 ( .A(n9068), .B(SI_26_), .ZN(n9070) );
  INV_X1 U10681 ( .A(n9070), .ZN(n9049) );
  XNOR2_X1 U10682 ( .A(n9071), .B(n9049), .ZN(n15122) );
  NAND2_X1 U10683 ( .A1(n15122), .A2(n9356), .ZN(n9051) );
  INV_X1 U10684 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n15125) );
  OR2_X1 U10685 ( .A1(n9357), .A2(n15125), .ZN(n9050) );
  XNOR2_X1 U10686 ( .A(n14856), .B(n14190), .ZN(n9064) );
  INV_X1 U10687 ( .A(n9054), .ZN(n9052) );
  INV_X1 U10688 ( .A(n9076), .ZN(n9078) );
  INV_X1 U10689 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9053) );
  NAND2_X1 U10690 ( .A1(n9054), .A2(n9053), .ZN(n9055) );
  NAND2_X1 U10691 ( .A1(n14854), .A2(n8836), .ZN(n9061) );
  INV_X1 U10692 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9058) );
  NAND2_X1 U10693 ( .A1(n9343), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U10694 ( .A1(n9342), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n9056) );
  OAI211_X1 U10695 ( .C1(n9058), .C2(n9346), .A(n9057), .B(n9056), .ZN(n9059)
         );
  INV_X1 U10696 ( .A(n9059), .ZN(n9060) );
  NAND2_X1 U10697 ( .A1(n14838), .A2(n14873), .ZN(n9065) );
  XNOR2_X1 U10698 ( .A(n9064), .B(n9065), .ZN(n14710) );
  AND2_X1 U10699 ( .A1(n14710), .A2(n9062), .ZN(n9063) );
  NAND2_X1 U10700 ( .A1(n14693), .A2(n9063), .ZN(n14699) );
  INV_X1 U10701 ( .A(n9064), .ZN(n9066) );
  NAND2_X1 U10702 ( .A1(n9066), .A2(n9065), .ZN(n9067) );
  NAND2_X1 U10703 ( .A1(n14699), .A2(n9067), .ZN(n9091) );
  NAND2_X1 U10704 ( .A1(n9068), .A2(SI_26_), .ZN(n9069) );
  INV_X1 U10705 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15980) );
  INV_X1 U10706 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n15120) );
  MUX2_X1 U10707 ( .A(n15980), .B(n15120), .S(n8511), .Z(n9296) );
  XNOR2_X1 U10708 ( .A(n9296), .B(SI_27_), .ZN(n9294) );
  INV_X1 U10709 ( .A(n9294), .ZN(n9072) );
  NAND2_X1 U10710 ( .A1(n15118), .A2(n9356), .ZN(n9074) );
  OR2_X1 U10711 ( .A1(n9357), .A2(n15120), .ZN(n9073) );
  XNOR2_X1 U10712 ( .A(n14843), .B(n9075), .ZN(n9086) );
  INV_X1 U10713 ( .A(n9138), .ZN(n9140) );
  INV_X1 U10714 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9077) );
  NAND2_X1 U10715 ( .A1(n9078), .A2(n9077), .ZN(n9079) );
  NAND2_X1 U10716 ( .A1(n14846), .A2(n8836), .ZN(n9085) );
  INV_X1 U10717 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9082) );
  NAND2_X1 U10718 ( .A1(n9343), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9081) );
  NAND2_X1 U10719 ( .A1(n9342), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9080) );
  OAI211_X1 U10720 ( .C1(n9082), .C2(n9346), .A(n9081), .B(n9080), .ZN(n9083)
         );
  INV_X1 U10721 ( .A(n9083), .ZN(n9084) );
  AND2_X1 U10722 ( .A1(n14861), .A2(n14986), .ZN(n9087) );
  NAND2_X1 U10723 ( .A1(n9086), .A2(n9087), .ZN(n14192) );
  INV_X1 U10724 ( .A(n9086), .ZN(n14187) );
  INV_X1 U10725 ( .A(n9087), .ZN(n9088) );
  NAND2_X1 U10726 ( .A1(n14187), .A2(n9088), .ZN(n9089) );
  NAND2_X1 U10727 ( .A1(n14192), .A2(n9089), .ZN(n9090) );
  OR2_X2 U10728 ( .A1(n9091), .A2(n9090), .ZN(n14193) );
  NAND2_X1 U10729 ( .A1(n9091), .A2(n9090), .ZN(n9128) );
  NOR4_X1 U10730 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n9100) );
  OR4_X1 U10731 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9097) );
  NOR4_X1 U10732 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n9095) );
  NOR4_X1 U10733 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9094) );
  NOR4_X1 U10734 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9093) );
  NOR4_X1 U10735 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9092) );
  NAND4_X1 U10736 ( .A1(n9095), .A2(n9094), .A3(n9093), .A4(n9092), .ZN(n9096)
         );
  NOR4_X1 U10737 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        n9097), .A4(n9096), .ZN(n9099) );
  NOR4_X1 U10738 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9098) );
  NAND3_X1 U10739 ( .A1(n9100), .A2(n9099), .A3(n9098), .ZN(n9115) );
  INV_X1 U10740 ( .A(n9101), .ZN(n9103) );
  NAND2_X1 U10741 ( .A1(n9112), .A2(n9111), .ZN(n9105) );
  OR2_X1 U10742 ( .A1(n9108), .A2(n9107), .ZN(n9109) );
  NAND2_X1 U10743 ( .A1(n9110), .A2(n9109), .ZN(n15127) );
  XNOR2_X1 U10744 ( .A(n15130), .B(P2_B_REG_SCAN_IN), .ZN(n9113) );
  NAND2_X1 U10745 ( .A1(n15127), .A2(n9113), .ZN(n9114) );
  AND2_X1 U10746 ( .A1(n9115), .A2(n16034), .ZN(n10446) );
  INV_X1 U10747 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n16038) );
  NAND2_X1 U10748 ( .A1(n16034), .A2(n16038), .ZN(n9118) );
  INV_X1 U10749 ( .A(n15130), .ZN(n9116) );
  OR2_X1 U10750 ( .A1(n15121), .A2(n9116), .ZN(n9117) );
  INV_X1 U10751 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n16033) );
  NAND2_X1 U10752 ( .A1(n16034), .A2(n16033), .ZN(n9121) );
  INV_X1 U10753 ( .A(n15127), .ZN(n9119) );
  OR2_X1 U10754 ( .A1(n15121), .A2(n9119), .ZN(n9120) );
  NAND2_X1 U10755 ( .A1(n9121), .A2(n9120), .ZN(n11315) );
  OR2_X1 U10756 ( .A1(n16039), .A2(n11315), .ZN(n9122) );
  NOR2_X1 U10757 ( .A1(n10446), .A2(n9122), .ZN(n9133) );
  NOR2_X1 U10758 ( .A1(n15127), .A2(n15130), .ZN(n9123) );
  NAND2_X1 U10759 ( .A1(n15121), .A2(n9123), .ZN(n10273) );
  NAND2_X1 U10760 ( .A1(n9124), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9126) );
  XNOR2_X1 U10761 ( .A(n9126), .B(n9125), .ZN(n9414) );
  NAND2_X1 U10762 ( .A1(n9155), .A2(n12727), .ZN(n9446) );
  NOR2_X1 U10763 ( .A1(n15079), .A2(n10269), .ZN(n9127) );
  INV_X1 U10764 ( .A(n14843), .ZN(n15016) );
  INV_X1 U10765 ( .A(n9129), .ZN(n9148) );
  NAND2_X1 U10766 ( .A1(n9130), .A2(n9441), .ZN(n11786) );
  OR2_X1 U10767 ( .A1(n9148), .A2(n11786), .ZN(n9132) );
  NAND2_X1 U10768 ( .A1(n14930), .A2(n11851), .ZN(n10447) );
  INV_X1 U10769 ( .A(n10447), .ZN(n9131) );
  INV_X1 U10770 ( .A(n9133), .ZN(n9134) );
  NAND2_X1 U10771 ( .A1(n9134), .A2(n10447), .ZN(n9137) );
  INV_X1 U10772 ( .A(n10445), .ZN(n9135) );
  AND2_X1 U10773 ( .A1(n10270), .A2(n9135), .ZN(n9136) );
  NAND2_X1 U10774 ( .A1(n9137), .A2(n9136), .ZN(n10661) );
  AOI22_X1 U10775 ( .A1(n14846), .A2(n14700), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9150) );
  NAND2_X1 U10776 ( .A1(n9138), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n12720) );
  INV_X1 U10777 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9139) );
  NAND2_X1 U10778 ( .A1(n9140), .A2(n9139), .ZN(n9141) );
  NAND2_X1 U10779 ( .A1(n12720), .A2(n9141), .ZN(n14194) );
  INV_X1 U10780 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9144) );
  NAND2_X1 U10781 ( .A1(n9343), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9143) );
  NAND2_X1 U10782 ( .A1(n9342), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9142) );
  OAI211_X1 U10783 ( .C1(n9144), .C2(n9346), .A(n9143), .B(n9142), .ZN(n9145)
         );
  INV_X1 U10784 ( .A(n9145), .ZN(n9146) );
  NAND2_X1 U10785 ( .A1(n10269), .A2(n15115), .ZN(n14953) );
  NOR2_X2 U10786 ( .A1(n14650), .A2(n14953), .ZN(n14702) );
  INV_X1 U10787 ( .A(n15115), .ZN(n10311) );
  NOR2_X2 U10788 ( .A1(n14650), .A2(n14951), .ZN(n14701) );
  AOI22_X1 U10789 ( .A1(n14839), .A2(n14702), .B1(n14701), .B2(n14838), .ZN(
        n9149) );
  OAI211_X1 U10790 ( .C1(n15016), .C2(n14705), .A(n9150), .B(n9149), .ZN(n9151) );
  INV_X1 U10791 ( .A(n9151), .ZN(n9152) );
  OAI21_X1 U10792 ( .B1(n14189), .B2(n9153), .A(n9152), .ZN(P2_U3186) );
  INV_X1 U10793 ( .A(n9156), .ZN(n9157) );
  NAND2_X1 U10794 ( .A1(n9370), .A2(n8032), .ZN(n9158) );
  INV_X1 U10795 ( .A(n11319), .ZN(n9403) );
  NAND2_X1 U10796 ( .A1(n14735), .A2(n9371), .ZN(n9165) );
  NAND2_X1 U10797 ( .A1(n9370), .A2(n16420), .ZN(n9164) );
  NAND2_X1 U10798 ( .A1(n14735), .A2(n9370), .ZN(n9167) );
  NAND2_X1 U10799 ( .A1(n9371), .A2(n16420), .ZN(n9166) );
  INV_X1 U10800 ( .A(n9222), .ZN(n9259) );
  NAND2_X1 U10801 ( .A1(n10716), .A2(n9259), .ZN(n9170) );
  NAND2_X1 U10802 ( .A1(n9170), .A2(n9169), .ZN(n9172) );
  AOI22_X1 U10804 ( .A1(n10716), .A2(n9222), .B1(n14734), .B2(n9259), .ZN(
        n9171) );
  INV_X1 U10805 ( .A(n9399), .ZN(n9372) );
  NAND2_X1 U10806 ( .A1(n14170), .A2(n9372), .ZN(n9175) );
  NAND2_X1 U10807 ( .A1(n14733), .A2(n9259), .ZN(n9174) );
  NAND2_X1 U10808 ( .A1(n9175), .A2(n9174), .ZN(n9177) );
  AOI22_X1 U10809 ( .A1(n14170), .A2(n9371), .B1(n9372), .B2(n14733), .ZN(
        n9176) );
  AOI21_X1 U10810 ( .B1(n9178), .B2(n9177), .A(n9176), .ZN(n9179) );
  NAND2_X1 U10811 ( .A1(n10998), .A2(n9259), .ZN(n9181) );
  NAND2_X1 U10812 ( .A1(n14732), .A2(n9361), .ZN(n9180) );
  AOI22_X1 U10813 ( .A1(n10998), .A2(n9361), .B1(n9371), .B2(n14732), .ZN(
        n9182) );
  NAND2_X1 U10814 ( .A1(n11802), .A2(n9361), .ZN(n9184) );
  NAND2_X1 U10815 ( .A1(n14731), .A2(n9259), .ZN(n9183) );
  NAND2_X1 U10816 ( .A1(n9184), .A2(n9183), .ZN(n9186) );
  AOI22_X1 U10817 ( .A1(n11802), .A2(n9371), .B1(n14731), .B2(n9361), .ZN(
        n9185) );
  AOI21_X1 U10818 ( .B1(n9187), .B2(n9186), .A(n9185), .ZN(n9189) );
  NOR2_X1 U10819 ( .A1(n9187), .A2(n9186), .ZN(n9188) );
  NAND2_X1 U10820 ( .A1(n11934), .A2(n9371), .ZN(n9191) );
  NAND2_X1 U10821 ( .A1(n14730), .A2(n9361), .ZN(n9190) );
  NAND2_X1 U10822 ( .A1(n9191), .A2(n9190), .ZN(n9194) );
  INV_X1 U10823 ( .A(n14730), .ZN(n11350) );
  NAND2_X1 U10824 ( .A1(n11934), .A2(n9361), .ZN(n9192) );
  OAI21_X1 U10825 ( .B1(n11350), .B2(n9370), .A(n9192), .ZN(n9193) );
  INV_X1 U10826 ( .A(n9194), .ZN(n9195) );
  NAND2_X1 U10827 ( .A1(n11548), .A2(n9361), .ZN(n9197) );
  NAND2_X1 U10828 ( .A1(n14729), .A2(n9259), .ZN(n9196) );
  NAND2_X1 U10829 ( .A1(n9197), .A2(n9196), .ZN(n9199) );
  AOI22_X1 U10830 ( .A1(n11548), .A2(n9371), .B1(n9361), .B2(n14729), .ZN(
        n9198) );
  NOR2_X1 U10831 ( .A1(n9200), .A2(n9199), .ZN(n9201) );
  OR2_X1 U10832 ( .A1(n9202), .A2(n9201), .ZN(n9207) );
  NAND2_X1 U10833 ( .A1(n12034), .A2(n9259), .ZN(n9204) );
  NAND2_X1 U10834 ( .A1(n14728), .A2(n9361), .ZN(n9203) );
  NAND2_X1 U10835 ( .A1(n9204), .A2(n9203), .ZN(n9208) );
  INV_X1 U10836 ( .A(n14728), .ZN(n11551) );
  NAND2_X1 U10837 ( .A1(n12034), .A2(n9361), .ZN(n9205) );
  OAI21_X1 U10838 ( .B1(n11551), .B2(n9370), .A(n9205), .ZN(n9206) );
  NAND2_X1 U10839 ( .A1(n12095), .A2(n9361), .ZN(n9210) );
  NAND2_X1 U10840 ( .A1(n14727), .A2(n9259), .ZN(n9209) );
  NAND2_X1 U10841 ( .A1(n9210), .A2(n9209), .ZN(n9212) );
  AOI22_X1 U10842 ( .A1(n12095), .A2(n9371), .B1(n9372), .B2(n14727), .ZN(
        n9211) );
  AOI21_X1 U10843 ( .B1(n9213), .B2(n9212), .A(n9211), .ZN(n9215) );
  NAND2_X1 U10844 ( .A1(n12151), .A2(n9259), .ZN(n9217) );
  NAND2_X1 U10845 ( .A1(n14726), .A2(n9361), .ZN(n9216) );
  NAND2_X1 U10846 ( .A1(n9217), .A2(n9216), .ZN(n9220) );
  AOI22_X1 U10847 ( .A1(n12151), .A2(n9361), .B1(n9371), .B2(n14726), .ZN(
        n9218) );
  INV_X1 U10848 ( .A(n9218), .ZN(n9219) );
  NAND2_X1 U10849 ( .A1(n12223), .A2(n9361), .ZN(n9224) );
  NAND2_X1 U10850 ( .A1(n14725), .A2(n9259), .ZN(n9223) );
  NAND2_X1 U10851 ( .A1(n9224), .A2(n9223), .ZN(n9227) );
  INV_X1 U10852 ( .A(n14725), .ZN(n11463) );
  NAND2_X1 U10853 ( .A1(n12223), .A2(n9399), .ZN(n9225) );
  OAI21_X1 U10854 ( .B1(n9399), .B2(n11463), .A(n9225), .ZN(n9226) );
  INV_X1 U10855 ( .A(n9226), .ZN(n9229) );
  NAND2_X1 U10856 ( .A1(n16606), .A2(n9259), .ZN(n9232) );
  NAND2_X1 U10857 ( .A1(n14724), .A2(n9361), .ZN(n9231) );
  NAND2_X1 U10858 ( .A1(n9232), .A2(n9231), .ZN(n9234) );
  AOI22_X1 U10859 ( .A1(n16606), .A2(n9361), .B1(n9371), .B2(n14724), .ZN(
        n9233) );
  NAND2_X1 U10860 ( .A1(n12427), .A2(n9361), .ZN(n9237) );
  NAND2_X1 U10861 ( .A1(n14723), .A2(n9399), .ZN(n9236) );
  NAND2_X1 U10862 ( .A1(n9237), .A2(n9236), .ZN(n9241) );
  INV_X1 U10863 ( .A(n14723), .ZN(n12369) );
  NAND2_X1 U10864 ( .A1(n12427), .A2(n9168), .ZN(n9238) );
  OAI21_X1 U10865 ( .B1(n9399), .B2(n12369), .A(n9238), .ZN(n9239) );
  NAND2_X1 U10866 ( .A1(n12566), .A2(n9399), .ZN(n9244) );
  NAND2_X1 U10867 ( .A1(n14722), .A2(n9361), .ZN(n9243) );
  AOI22_X1 U10868 ( .A1(n12566), .A2(n9361), .B1(n9371), .B2(n14722), .ZN(
        n9245) );
  NAND2_X1 U10869 ( .A1(n15078), .A2(n9361), .ZN(n9247) );
  NAND2_X1 U10870 ( .A1(n14721), .A2(n9371), .ZN(n9246) );
  NAND2_X1 U10871 ( .A1(n9247), .A2(n9246), .ZN(n9250) );
  INV_X1 U10872 ( .A(n14721), .ZN(n12626) );
  NAND2_X1 U10873 ( .A1(n15078), .A2(n9259), .ZN(n9248) );
  OAI21_X1 U10874 ( .B1(n9399), .B2(n12626), .A(n9248), .ZN(n9249) );
  NAND2_X1 U10875 ( .A1(n15073), .A2(n9259), .ZN(n9252) );
  NAND2_X1 U10876 ( .A1(n14720), .A2(n9222), .ZN(n9251) );
  AOI22_X1 U10877 ( .A1(n15073), .A2(n9361), .B1(n9371), .B2(n14720), .ZN(
        n9253) );
  NAND2_X1 U10878 ( .A1(n15068), .A2(n9361), .ZN(n9255) );
  NAND2_X1 U10879 ( .A1(n14719), .A2(n9168), .ZN(n9254) );
  NAND2_X1 U10880 ( .A1(n9255), .A2(n9254), .ZN(n9257) );
  AOI22_X1 U10881 ( .A1(n15068), .A2(n9371), .B1(n9370), .B2(n14719), .ZN(
        n9256) );
  NAND2_X1 U10882 ( .A1(n15062), .A2(n9259), .ZN(n9261) );
  NAND2_X1 U10883 ( .A1(n14718), .A2(n9361), .ZN(n9260) );
  NAND2_X1 U10884 ( .A1(n9261), .A2(n9260), .ZN(n9264) );
  NAND2_X1 U10885 ( .A1(n15062), .A2(n9372), .ZN(n9262) );
  OAI21_X1 U10886 ( .B1(n14177), .B2(n9370), .A(n9262), .ZN(n9263) );
  NAND2_X1 U10887 ( .A1(n15057), .A2(n9372), .ZN(n9267) );
  NAND2_X1 U10888 ( .A1(n14717), .A2(n9371), .ZN(n9266) );
  NAND2_X1 U10889 ( .A1(n9267), .A2(n9266), .ZN(n9269) );
  AOI22_X1 U10890 ( .A1(n15057), .A2(n9371), .B1(n9370), .B2(n14717), .ZN(
        n9268) );
  INV_X1 U10891 ( .A(n9274), .ZN(n9271) );
  AND2_X1 U10892 ( .A1(n14716), .A2(n9361), .ZN(n9270) );
  AOI21_X1 U10893 ( .B1(n15053), .B2(n9371), .A(n9270), .ZN(n9272) );
  NAND2_X1 U10894 ( .A1(n9271), .A2(n9272), .ZN(n9280) );
  INV_X1 U10895 ( .A(n9272), .ZN(n9273) );
  NAND2_X1 U10896 ( .A1(n9274), .A2(n9273), .ZN(n9278) );
  NAND2_X1 U10897 ( .A1(n15053), .A2(n9361), .ZN(n9276) );
  NAND2_X1 U10898 ( .A1(n14716), .A2(n9371), .ZN(n9275) );
  NAND2_X1 U10899 ( .A1(n9276), .A2(n9275), .ZN(n9277) );
  NAND2_X1 U10900 ( .A1(n9278), .A2(n9277), .ZN(n9279) );
  NAND2_X1 U10901 ( .A1(n15048), .A2(n9372), .ZN(n9282) );
  NAND2_X1 U10902 ( .A1(n14912), .A2(n9371), .ZN(n9281) );
  NAND2_X1 U10903 ( .A1(n9282), .A2(n9281), .ZN(n9284) );
  AOI22_X1 U10904 ( .A1(n15048), .A2(n9371), .B1(n9361), .B2(n14912), .ZN(
        n9283) );
  NAND2_X1 U10905 ( .A1(n15039), .A2(n9371), .ZN(n9286) );
  NAND2_X1 U10906 ( .A1(n14715), .A2(n9370), .ZN(n9285) );
  AOI22_X1 U10907 ( .A1(n15039), .A2(n9361), .B1(n9371), .B2(n14715), .ZN(
        n9287) );
  AOI22_X1 U10908 ( .A1(n15035), .A2(n9361), .B1(n9371), .B2(n14914), .ZN(
        n9289) );
  AOI22_X1 U10909 ( .A1(n15035), .A2(n9371), .B1(n9361), .B2(n14914), .ZN(
        n9291) );
  OAI22_X1 U10910 ( .A1(n14889), .A2(n9370), .B1(n9399), .B2(n14870), .ZN(
        n9293) );
  AOI22_X1 U10911 ( .A1(n7953), .A2(n9361), .B1(n9371), .B2(n14860), .ZN(n9374) );
  OAI22_X1 U10912 ( .A1(n14877), .A2(n9370), .B1(n9399), .B2(n14695), .ZN(
        n9373) );
  AOI22_X1 U10913 ( .A1(n15030), .A2(n9370), .B1(n9371), .B2(n14714), .ZN(
        n9292) );
  INV_X1 U10914 ( .A(n9296), .ZN(n9297) );
  INV_X1 U10915 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13372) );
  INV_X1 U10916 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n15117) );
  MUX2_X1 U10917 ( .A(n13372), .B(n15117), .S(n8511), .Z(n9298) );
  INV_X1 U10918 ( .A(SI_28_), .ZN(n14407) );
  NAND2_X1 U10919 ( .A1(n9298), .A2(n14407), .ZN(n9301) );
  INV_X1 U10920 ( .A(n9298), .ZN(n9299) );
  NAND2_X1 U10921 ( .A1(n9299), .A2(SI_28_), .ZN(n9300) );
  NAND2_X1 U10922 ( .A1(n9301), .A2(n9300), .ZN(n9354) );
  INV_X1 U10923 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15977) );
  INV_X1 U10924 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n15113) );
  MUX2_X1 U10925 ( .A(n15977), .B(n15113), .S(n8511), .Z(n9302) );
  XNOR2_X1 U10926 ( .A(n9302), .B(SI_29_), .ZN(n9337) );
  INV_X1 U10927 ( .A(n9302), .ZN(n9303) );
  NOR2_X1 U10928 ( .A1(n9303), .A2(SI_29_), .ZN(n9304) );
  MUX2_X1 U10929 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8511), .Z(n9305) );
  NAND2_X1 U10930 ( .A1(n9305), .A2(SI_30_), .ZN(n9307) );
  OAI21_X1 U10931 ( .B1(n9305), .B2(SI_30_), .A(n9307), .ZN(n9317) );
  INV_X1 U10932 ( .A(n9317), .ZN(n9306) );
  NAND2_X1 U10933 ( .A1(n9316), .A2(n9306), .ZN(n9320) );
  NAND2_X1 U10934 ( .A1(n9320), .A2(n9307), .ZN(n9310) );
  MUX2_X1 U10935 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10468), .Z(n9308) );
  XNOR2_X1 U10936 ( .A(n9308), .B(SI_31_), .ZN(n9309) );
  NAND2_X1 U10937 ( .A1(n15104), .A2(n9356), .ZN(n9312) );
  INV_X1 U10938 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n15107) );
  OR2_X1 U10939 ( .A1(n9357), .A2(n15107), .ZN(n9311) );
  INV_X1 U10940 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9315) );
  NAND2_X1 U10941 ( .A1(n9343), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9314) );
  NAND2_X1 U10942 ( .A1(n9342), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9313) );
  OAI211_X1 U10943 ( .C1(n9346), .C2(n9315), .A(n9314), .B(n9313), .ZN(n14807)
         );
  INV_X1 U10944 ( .A(n9316), .ZN(n9318) );
  NAND2_X1 U10945 ( .A1(n9318), .A2(n9317), .ZN(n9319) );
  INV_X1 U10946 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12731) );
  OR2_X1 U10947 ( .A1(n9357), .A2(n12731), .ZN(n9322) );
  NAND2_X1 U10948 ( .A1(n14807), .A2(n9372), .ZN(n9398) );
  AND2_X1 U10949 ( .A1(n9446), .A2(n9405), .ZN(n9324) );
  OR2_X1 U10950 ( .A1(n11323), .A2(n9157), .ZN(n9408) );
  AND2_X1 U10951 ( .A1(n9324), .A2(n9408), .ZN(n9332) );
  INV_X1 U10952 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9325) );
  OR2_X1 U10953 ( .A1(n8620), .A2(n9325), .ZN(n9331) );
  INV_X1 U10954 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n9326) );
  OR2_X1 U10955 ( .A1(n9327), .A2(n9326), .ZN(n9330) );
  INV_X1 U10956 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9328) );
  OR2_X1 U10957 ( .A1(n9346), .A2(n9328), .ZN(n9329) );
  AND3_X1 U10958 ( .A1(n9331), .A2(n9330), .A3(n9329), .ZN(n9334) );
  AOI21_X1 U10959 ( .B1(n9398), .B2(n9332), .A(n9334), .ZN(n9333) );
  AOI21_X1 U10960 ( .B1(n14810), .B2(n9371), .A(n9333), .ZN(n9391) );
  NAND2_X1 U10961 ( .A1(n14810), .A2(n9372), .ZN(n9336) );
  INV_X1 U10962 ( .A(n9334), .ZN(n14712) );
  NAND2_X1 U10963 ( .A1(n14712), .A2(n9259), .ZN(n9335) );
  NAND2_X1 U10964 ( .A1(n9336), .A2(n9335), .ZN(n9390) );
  NAND2_X1 U10965 ( .A1(n15112), .A2(n9356), .ZN(n9340) );
  OR2_X1 U10966 ( .A1(n9357), .A2(n15113), .ZN(n9339) );
  OR2_X1 U10967 ( .A1(n12720), .A2(n9341), .ZN(n9350) );
  INV_X1 U10968 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9347) );
  NAND2_X1 U10969 ( .A1(n9342), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n9345) );
  NAND2_X1 U10970 ( .A1(n9343), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9344) );
  OAI211_X1 U10971 ( .C1(n9347), .C2(n9346), .A(n9345), .B(n9344), .ZN(n9348)
         );
  INV_X1 U10972 ( .A(n9348), .ZN(n9349) );
  NAND2_X1 U10973 ( .A1(n9350), .A2(n9349), .ZN(n14713) );
  AND2_X1 U10974 ( .A1(n14713), .A2(n9372), .ZN(n9351) );
  AOI21_X1 U10975 ( .B1(n15005), .B2(n9371), .A(n9351), .ZN(n9382) );
  NAND2_X1 U10976 ( .A1(n15005), .A2(n9361), .ZN(n9353) );
  NAND2_X1 U10977 ( .A1(n14713), .A2(n9371), .ZN(n9352) );
  NAND2_X1 U10978 ( .A1(n9353), .A2(n9352), .ZN(n9381) );
  NAND2_X1 U10979 ( .A1(n13371), .A2(n9356), .ZN(n9359) );
  OR2_X1 U10980 ( .A1(n9357), .A2(n15117), .ZN(n9358) );
  AND2_X1 U10981 ( .A1(n14839), .A2(n9371), .ZN(n9360) );
  AOI21_X1 U10982 ( .B1(n15011), .B2(n9361), .A(n9360), .ZN(n9378) );
  NAND2_X1 U10983 ( .A1(n15011), .A2(n9371), .ZN(n9363) );
  NAND2_X1 U10984 ( .A1(n14839), .A2(n9222), .ZN(n9362) );
  NAND2_X1 U10985 ( .A1(n9363), .A2(n9362), .ZN(n9377) );
  NAND2_X1 U10986 ( .A1(n9378), .A2(n9377), .ZN(n9364) );
  NAND2_X1 U10987 ( .A1(n9383), .A2(n9364), .ZN(n9388) );
  AND2_X1 U10988 ( .A1(n14861), .A2(n9371), .ZN(n9365) );
  AOI21_X1 U10989 ( .B1(n14843), .B2(n9372), .A(n9365), .ZN(n9387) );
  NAND2_X1 U10990 ( .A1(n14843), .A2(n9371), .ZN(n9368) );
  NAND2_X1 U10991 ( .A1(n14861), .A2(n9372), .ZN(n9367) );
  NAND2_X1 U10992 ( .A1(n9368), .A2(n9367), .ZN(n9386) );
  AND2_X1 U10993 ( .A1(n9387), .A2(n9386), .ZN(n9369) );
  OAI22_X1 U10994 ( .A1(n14856), .A2(n9370), .B1(n9399), .B2(n14871), .ZN(
        n9392) );
  AOI22_X1 U10995 ( .A1(n15022), .A2(n9372), .B1(n9371), .B2(n14838), .ZN(
        n9393) );
  AOI22_X1 U10996 ( .A1(n9392), .A2(n9393), .B1(n9374), .B2(n9373), .ZN(n9375)
         );
  INV_X1 U10997 ( .A(n9377), .ZN(n9380) );
  INV_X1 U10998 ( .A(n9378), .ZN(n9379) );
  AOI22_X1 U10999 ( .A1(n9382), .A2(n9381), .B1(n9380), .B2(n9379), .ZN(n9385)
         );
  INV_X1 U11000 ( .A(n9383), .ZN(n9384) );
  AOI21_X1 U11001 ( .B1(n9385), .B2(n9415), .A(n9384), .ZN(n9389) );
  INV_X1 U11002 ( .A(n9392), .ZN(n9395) );
  INV_X1 U11003 ( .A(n9393), .ZN(n9394) );
  NAND3_X1 U11004 ( .A1(n9396), .A2(n9395), .A3(n9394), .ZN(n9397) );
  NAND2_X1 U11005 ( .A1(n9398), .A2(n9361), .ZN(n9401) );
  NAND2_X1 U11006 ( .A1(n9399), .A2(n14807), .ZN(n9400) );
  MUX2_X1 U11007 ( .A(n9401), .B(n9400), .S(n15000), .Z(n9402) );
  OAI21_X1 U11008 ( .B1(n9403), .B2(n8519), .A(n11851), .ZN(n9404) );
  OAI21_X1 U11009 ( .B1(n9155), .B2(n9405), .A(n9404), .ZN(n9406) );
  INV_X1 U11010 ( .A(n9408), .ZN(n9410) );
  NOR3_X1 U11011 ( .A1(n9155), .A2(n12139), .A3(n12727), .ZN(n9409) );
  NOR2_X1 U11012 ( .A1(n9410), .A2(n9409), .ZN(n9411) );
  INV_X1 U11013 ( .A(n9414), .ZN(n10272) );
  AND2_X1 U11014 ( .A1(n10272), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9439) );
  INV_X1 U11015 ( .A(n9439), .ZN(n12471) );
  INV_X1 U11016 ( .A(n9415), .ZN(n9438) );
  INV_X1 U11017 ( .A(n14713), .ZN(n14820) );
  XNOR2_X1 U11018 ( .A(n15005), .B(n14820), .ZN(n12716) );
  XNOR2_X1 U11019 ( .A(n14810), .B(n14712), .ZN(n9436) );
  INV_X1 U11020 ( .A(n14839), .ZN(n9416) );
  NAND2_X1 U11021 ( .A1(n15011), .A2(n9416), .ZN(n9417) );
  NAND2_X1 U11022 ( .A1(n15022), .A2(n14871), .ZN(n12689) );
  OR2_X1 U11023 ( .A1(n15022), .A2(n14871), .ZN(n9418) );
  NAND2_X1 U11024 ( .A1(n12689), .A2(n9418), .ZN(n12688) );
  NAND2_X1 U11025 ( .A1(n7953), .A2(n14860), .ZN(n12710) );
  NAND2_X1 U11026 ( .A1(n12711), .A2(n12710), .ZN(n14868) );
  XNOR2_X1 U11027 ( .A(n15039), .B(n14942), .ZN(n12706) );
  XNOR2_X1 U11028 ( .A(n15048), .B(n14912), .ZN(n14938) );
  XNOR2_X1 U11029 ( .A(n15062), .B(n14177), .ZN(n14984) );
  XNOR2_X1 U11030 ( .A(n15068), .B(n14719), .ZN(n12642) );
  XNOR2_X1 U11031 ( .A(n12566), .B(n12571), .ZN(n12376) );
  XNOR2_X1 U11032 ( .A(n12427), .B(n14723), .ZN(n12267) );
  INV_X1 U11033 ( .A(n14724), .ZN(n12265) );
  NAND2_X1 U11034 ( .A1(n16606), .A2(n12265), .ZN(n12268) );
  OR2_X1 U11035 ( .A1(n16606), .A2(n12265), .ZN(n9419) );
  NAND2_X1 U11036 ( .A1(n12223), .A2(n11463), .ZN(n12191) );
  OR2_X1 U11037 ( .A1(n12223), .A2(n11463), .ZN(n9420) );
  NAND2_X1 U11038 ( .A1(n12191), .A2(n9420), .ZN(n12073) );
  XNOR2_X1 U11039 ( .A(n12034), .B(n14728), .ZN(n12033) );
  INV_X1 U11040 ( .A(n14737), .ZN(n10625) );
  NAND2_X1 U11041 ( .A1(n10625), .A2(n8032), .ZN(n10659) );
  AND2_X1 U11042 ( .A1(n9421), .A2(n10659), .ZN(n11328) );
  NAND4_X1 U11043 ( .A1(n11328), .A2(n9441), .A3(n10610), .A4(n10622), .ZN(
        n9423) );
  XNOR2_X1 U11044 ( .A(n11802), .B(n14731), .ZN(n11000) );
  NAND2_X1 U11045 ( .A1(n10815), .A2(n11000), .ZN(n9422) );
  NOR2_X1 U11046 ( .A1(n9423), .A2(n9422), .ZN(n9424) );
  XNOR2_X1 U11047 ( .A(n10998), .B(n14732), .ZN(n10995) );
  NAND4_X1 U11048 ( .A1(n12033), .A2(n9424), .A3(n10995), .A4(n11918), .ZN(
        n9425) );
  XNOR2_X1 U11049 ( .A(n12095), .B(n12065), .ZN(n12069) );
  XNOR2_X1 U11050 ( .A(n11548), .B(n12029), .ZN(n11353) );
  OR3_X1 U11051 ( .A1(n9425), .A2(n12069), .A3(n11353), .ZN(n9426) );
  NOR2_X1 U11052 ( .A1(n12073), .A2(n9426), .ZN(n9427) );
  XNOR2_X1 U11053 ( .A(n12151), .B(n14726), .ZN(n12144) );
  NAND4_X1 U11054 ( .A1(n12267), .A2(n12194), .A3(n9427), .A4(n12144), .ZN(
        n9428) );
  NOR2_X1 U11055 ( .A1(n12376), .A2(n9428), .ZN(n9429) );
  XNOR2_X1 U11056 ( .A(n15073), .B(n14720), .ZN(n12594) );
  XNOR2_X1 U11057 ( .A(n15078), .B(n14721), .ZN(n12569) );
  NAND4_X1 U11058 ( .A1(n12642), .A2(n9429), .A3(n12594), .A4(n12569), .ZN(
        n9430) );
  NOR2_X1 U11059 ( .A1(n14984), .A2(n9430), .ZN(n9431) );
  XNOR2_X1 U11060 ( .A(n15053), .B(n14716), .ZN(n14947) );
  XNOR2_X1 U11061 ( .A(n15057), .B(n14717), .ZN(n14967) );
  NAND4_X1 U11062 ( .A1(n14938), .A2(n9431), .A3(n14947), .A4(n14967), .ZN(
        n9432) );
  NOR2_X1 U11063 ( .A1(n12706), .A2(n9432), .ZN(n9433) );
  XNOR2_X1 U11064 ( .A(n15030), .B(n14714), .ZN(n14891) );
  XNOR2_X1 U11065 ( .A(n15035), .B(n14914), .ZN(n14900) );
  NAND4_X1 U11066 ( .A1(n14868), .A2(n9433), .A3(n14891), .A4(n14900), .ZN(
        n9434) );
  NOR2_X1 U11067 ( .A1(n12688), .A2(n9434), .ZN(n9435) );
  NAND4_X1 U11068 ( .A1(n9436), .A2(n14822), .A3(n9435), .A4(n14834), .ZN(
        n9437) );
  NOR3_X1 U11069 ( .A1(n9438), .A2(n12716), .A3(n9437), .ZN(n9445) );
  NAND2_X1 U11070 ( .A1(n9439), .A2(n12139), .ZN(n9443) );
  NOR3_X1 U11071 ( .A1(n9445), .A2(n12727), .A3(n9443), .ZN(n9440) );
  OAI21_X1 U11072 ( .B1(n9442), .B2(n9441), .A(n9440), .ZN(n9452) );
  INV_X1 U11073 ( .A(n9443), .ZN(n9444) );
  INV_X1 U11074 ( .A(n9446), .ZN(n9447) );
  INV_X1 U11075 ( .A(n15119), .ZN(n10306) );
  NAND4_X1 U11076 ( .A1(n16040), .A2(n9447), .A3(n10306), .A4(n14911), .ZN(
        n9448) );
  OAI211_X1 U11077 ( .C1(n8519), .C2(n12471), .A(n9448), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9449) );
  INV_X1 U11078 ( .A(n9449), .ZN(n9450) );
  AND2_X1 U11079 ( .A1(n9452), .A2(n9451), .ZN(n9453) );
  OAI21_X1 U11080 ( .B1(n9454), .B2(n12471), .A(n9453), .ZN(P2_U3328) );
  INV_X1 U11081 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n10087) );
  INV_X1 U11082 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n9616) );
  NAND2_X1 U11083 ( .A1(n9460), .A2(n9459), .ZN(n9765) );
  INV_X1 U11084 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9461) );
  NAND2_X1 U11085 ( .A1(n9807), .A2(n9461), .ZN(n9824) );
  INV_X1 U11086 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n9462) );
  INV_X1 U11087 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9463) );
  NOR2_X1 U11088 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), 
        .ZN(n9467) );
  NOR2_X1 U11089 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), 
        .ZN(n9466) );
  NOR2_X1 U11090 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), 
        .ZN(n9465) );
  NAND2_X1 U11091 ( .A1(n9464), .A2(n9547), .ZN(n9469) );
  NAND2_X1 U11092 ( .A1(n9469), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9468) );
  MUX2_X1 U11093 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9468), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n9471) );
  INV_X1 U11094 ( .A(n9469), .ZN(n9470) );
  NAND2_X1 U11095 ( .A1(n9471), .A2(n9473), .ZN(n11281) );
  NAND2_X1 U11096 ( .A1(n13694), .A2(n11281), .ZN(n10094) );
  NAND2_X1 U11097 ( .A1(n10074), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9472) );
  NAND2_X1 U11098 ( .A1(n13706), .A2(n12963), .ZN(n10096) );
  NAND2_X1 U11099 ( .A1(n10094), .A2(n10096), .ZN(n10082) );
  OR2_X1 U11100 ( .A1(n10082), .A2(n9480), .ZN(n10050) );
  NAND2_X1 U11101 ( .A1(n9473), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9474) );
  MUX2_X1 U11102 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9474), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n9475) );
  NAND2_X1 U11103 ( .A1(n13694), .A2(n11442), .ZN(n9478) );
  AND2_X1 U11104 ( .A1(n11442), .A2(n11281), .ZN(n10084) );
  INV_X1 U11105 ( .A(n10084), .ZN(n9476) );
  XNOR2_X1 U11106 ( .A(n12963), .B(n9476), .ZN(n9477) );
  NAND2_X1 U11107 ( .A1(n9478), .A2(n9477), .ZN(n10728) );
  INV_X1 U11108 ( .A(n10094), .ZN(n12921) );
  NAND3_X1 U11109 ( .A1(n10728), .A2(n12921), .A3(n16580), .ZN(n9479) );
  AND2_X1 U11110 ( .A1(n12920), .A2(n9480), .ZN(n16485) );
  XNOR2_X1 U11111 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9602) );
  AND2_X2 U11112 ( .A1(n9481), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9601) );
  NAND2_X1 U11113 ( .A1(n9602), .A2(n9601), .ZN(n9483) );
  NAND2_X1 U11114 ( .A1(n10146), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9482) );
  NAND2_X1 U11115 ( .A1(n10172), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9486) );
  NAND2_X1 U11116 ( .A1(n10493), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n9484) );
  NAND2_X1 U11117 ( .A1(n9486), .A2(n9484), .ZN(n9612) );
  INV_X1 U11118 ( .A(n9612), .ZN(n9485) );
  NAND2_X1 U11119 ( .A1(n9613), .A2(n9485), .ZN(n9487) );
  NAND2_X1 U11120 ( .A1(n9487), .A2(n9486), .ZN(n9623) );
  NAND2_X1 U11121 ( .A1(n10164), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9489) );
  NAND2_X1 U11122 ( .A1(n7671), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n9488) );
  NAND2_X1 U11123 ( .A1(n9623), .A2(n9622), .ZN(n9490) );
  NAND2_X1 U11124 ( .A1(n10186), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n9491) );
  NAND2_X1 U11125 ( .A1(n9638), .A2(n9637), .ZN(n9493) );
  NAND2_X1 U11126 ( .A1(n10195), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n9494) );
  NAND2_X1 U11127 ( .A1(n9496), .A2(n9494), .ZN(n9655) );
  INV_X1 U11128 ( .A(n9655), .ZN(n9495) );
  NAND2_X1 U11129 ( .A1(n9656), .A2(n9495), .ZN(n9497) );
  NAND2_X1 U11130 ( .A1(n10192), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9498) );
  NAND2_X1 U11131 ( .A1(n9670), .A2(n9498), .ZN(n9500) );
  NAND2_X1 U11132 ( .A1(n10173), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9499) );
  NAND2_X1 U11133 ( .A1(n10209), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n9501) );
  NAND2_X1 U11134 ( .A1(n9502), .A2(n9501), .ZN(n9681) );
  NAND2_X1 U11135 ( .A1(n9504), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n9505) );
  NAND2_X1 U11136 ( .A1(n10229), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n9506) );
  NAND2_X1 U11137 ( .A1(n9507), .A2(n9506), .ZN(n9711) );
  NAND2_X1 U11138 ( .A1(n10235), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9509) );
  NAND2_X1 U11139 ( .A1(n10231), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n9508) );
  XNOR2_X1 U11140 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9745) );
  INV_X1 U11141 ( .A(n9745), .ZN(n9510) );
  INV_X1 U11142 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U11143 ( .A1(n9511), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n9512) );
  NAND2_X1 U11144 ( .A1(n10252), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9514) );
  NAND2_X1 U11145 ( .A1(n10248), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n9513) );
  XNOR2_X1 U11146 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n9790) );
  INV_X1 U11147 ( .A(n9790), .ZN(n9515) );
  NAND2_X1 U11148 ( .A1(n10650), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9517) );
  NAND2_X1 U11149 ( .A1(n10643), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n9516) );
  NAND2_X1 U11150 ( .A1(n9517), .A2(n9516), .ZN(n9803) );
  OR2_X2 U11151 ( .A1(n9804), .A2(n9803), .ZN(n9806) );
  NAND2_X1 U11152 ( .A1(n11012), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9520) );
  NAND2_X1 U11153 ( .A1(n10889), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n9518) );
  NAND2_X1 U11154 ( .A1(n9520), .A2(n9518), .ZN(n9820) );
  INV_X1 U11155 ( .A(n9820), .ZN(n9519) );
  NAND2_X2 U11156 ( .A1(n9819), .A2(n9519), .ZN(n9822) );
  INV_X1 U11157 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9521) );
  XNOR2_X1 U11158 ( .A(n9521), .B(P2_DATAO_REG_17__SCAN_IN), .ZN(n9838) );
  NAND2_X1 U11159 ( .A1(n11473), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9523) );
  NAND2_X1 U11160 ( .A1(n11495), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n9522) );
  NAND2_X1 U11161 ( .A1(n9523), .A2(n9522), .ZN(n9853) );
  INV_X1 U11162 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11701) );
  NAND2_X1 U11163 ( .A1(n11701), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9525) );
  INV_X1 U11164 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12729) );
  NAND2_X1 U11165 ( .A1(n12729), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9524) );
  XNOR2_X1 U11166 ( .A(n12045), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n9882) );
  NAND2_X1 U11167 ( .A1(n12045), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9526) );
  INV_X1 U11168 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n13183) );
  NAND2_X1 U11169 ( .A1(n13183), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9528) );
  NAND2_X1 U11170 ( .A1(n12141), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9527) );
  AND2_X1 U11171 ( .A1(n9528), .A2(n9527), .ZN(n9893) );
  INV_X1 U11172 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9529) );
  NAND2_X1 U11173 ( .A1(n9529), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9532) );
  NAND2_X1 U11174 ( .A1(n12298), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9530) );
  NAND2_X1 U11175 ( .A1(n9532), .A2(n9530), .ZN(n9905) );
  INV_X1 U11176 ( .A(n9905), .ZN(n9531) );
  NAND2_X1 U11177 ( .A1(n9906), .A2(n9531), .ZN(n9533) );
  XNOR2_X1 U11178 ( .A(n12473), .B(P2_DATAO_REG_23__SCAN_IN), .ZN(n9916) );
  NAND2_X1 U11179 ( .A1(n12473), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9534) );
  INV_X1 U11180 ( .A(n9925), .ZN(n9537) );
  NOR2_X2 U11181 ( .A1(n9535), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9536) );
  NAND2_X1 U11182 ( .A1(n15988), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9540) );
  NAND2_X1 U11183 ( .A1(n15128), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9538) );
  NAND2_X1 U11184 ( .A1(n9540), .A2(n9538), .ZN(n9933) );
  INV_X1 U11185 ( .A(n9933), .ZN(n9539) );
  INV_X1 U11186 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15983) );
  NAND2_X1 U11187 ( .A1(n15983), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9542) );
  NAND2_X1 U11188 ( .A1(n15125), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9541) );
  AND2_X1 U11189 ( .A1(n9542), .A2(n9541), .ZN(n9947) );
  NAND2_X1 U11190 ( .A1(n15980), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9544) );
  NAND2_X1 U11191 ( .A1(n15120), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9543) );
  AND2_X1 U11192 ( .A1(n9544), .A2(n9543), .ZN(n9961) );
  NAND2_X1 U11193 ( .A1(n13372), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9546) );
  NAND2_X1 U11194 ( .A1(n15117), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9545) );
  AND2_X1 U11195 ( .A1(n9546), .A2(n9545), .ZN(n9976) );
  XNOR2_X1 U11196 ( .A(n15977), .B(P1_DATAO_REG_29__SCAN_IN), .ZN(n12744) );
  XNOR2_X1 U11197 ( .A(n12746), .B(n12744), .ZN(n14149) );
  NAND4_X1 U11198 ( .A1(n9548), .A2(n9549), .A3(n9550), .A4(n10075), .ZN(n9551) );
  XNOR2_X2 U11199 ( .A(n9557), .B(n9556), .ZN(n10036) );
  NAND2_X1 U11200 ( .A1(n14149), .A2(n12759), .ZN(n9559) );
  NAND2_X1 U11201 ( .A1(n12760), .A2(SI_29_), .ZN(n9558) );
  NAND2_X1 U11202 ( .A1(n9559), .A2(n9558), .ZN(n10088) );
  NOR2_X1 U11203 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_REG3_REG_5__SCAN_IN), 
        .ZN(n9560) );
  NAND2_X1 U11204 ( .A1(n9561), .A2(n9560), .ZN(n9675) );
  INV_X1 U11205 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n13511) );
  INV_X1 U11206 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n14295) );
  INV_X1 U11207 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n14291) );
  INV_X1 U11208 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n14497) );
  INV_X1 U11209 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9570) );
  INV_X1 U11210 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n14505) );
  INV_X1 U11211 ( .A(n9982), .ZN(n9573) );
  INV_X1 U11212 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n13430) );
  NAND2_X1 U11213 ( .A1(n9573), .A2(n13430), .ZN(n13718) );
  OR2_X2 U11214 ( .A1(n9577), .A2(n14143), .ZN(n9574) );
  XNOR2_X2 U11215 ( .A(n9574), .B(P3_IR_REG_30__SCAN_IN), .ZN(n9579) );
  INV_X1 U11216 ( .A(n9577), .ZN(n14144) );
  OR2_X1 U11217 ( .A1(n13718), .A2(n9662), .ZN(n12743) );
  INV_X1 U11218 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n9583) );
  NAND2_X1 U11219 ( .A1(n10038), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9582) );
  NAND2_X1 U11220 ( .A1(n9954), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9581) );
  OAI211_X1 U11221 ( .C1(n9583), .C2(n7436), .A(n9582), .B(n9581), .ZN(n9584)
         );
  INV_X1 U11222 ( .A(n9584), .ZN(n9585) );
  OR2_X2 U11223 ( .A1(n10088), .A2(n13734), .ZN(n12904) );
  NAND2_X1 U11224 ( .A1(n10088), .A2(n13734), .ZN(n12906) );
  NAND2_X1 U11225 ( .A1(n10039), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9589) );
  NAND2_X1 U11226 ( .A1(n7437), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9588) );
  INV_X1 U11227 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9586) );
  NAND2_X1 U11228 ( .A1(n7435), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9590) );
  INV_X1 U11229 ( .A(n10636), .ZN(n9598) );
  INV_X1 U11230 ( .A(n9644), .ZN(n9595) );
  INV_X1 U11231 ( .A(n9601), .ZN(n9594) );
  NAND2_X1 U11232 ( .A1(n9592), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9593) );
  NAND2_X1 U11233 ( .A1(n9594), .A2(n9593), .ZN(n10156) );
  NAND2_X1 U11234 ( .A1(n9595), .A2(n10156), .ZN(n9597) );
  NAND2_X1 U11235 ( .A1(n9768), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U11236 ( .A1(n9984), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9606) );
  NAND2_X1 U11237 ( .A1(n7437), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n9605) );
  INV_X1 U11238 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n9599) );
  INV_X1 U11239 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11536) );
  NAND2_X1 U11240 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n9600) );
  XNOR2_X1 U11241 ( .A(n9602), .B(n9601), .ZN(n9603) );
  MUX2_X1 U11242 ( .A(n9603), .B(SI_1_), .S(n10468), .Z(n14156) );
  MUX2_X1 U11243 ( .A(n14155), .B(n14156), .S(n10928), .Z(n11033) );
  NAND2_X1 U11244 ( .A1(n11537), .A2(n9990), .ZN(n9607) );
  NAND4_X1 U11245 ( .A1(n9606), .A2(n9605), .A3(n9604), .A4(n7443), .ZN(n10734) );
  INV_X1 U11246 ( .A(n11033), .ZN(n11529) );
  NAND2_X1 U11247 ( .A1(n10734), .A2(n11529), .ZN(n12788) );
  NAND2_X1 U11248 ( .A1(n10038), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9611) );
  INV_X1 U11249 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10932) );
  OR2_X1 U11250 ( .A1(n7436), .A2(n10932), .ZN(n9610) );
  NAND2_X1 U11251 ( .A1(n10039), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n9609) );
  NAND2_X1 U11252 ( .A1(n7437), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n9608) );
  XNOR2_X1 U11253 ( .A(n9612), .B(n9613), .ZN(n10149) );
  INV_X1 U11254 ( .A(n10149), .ZN(n9614) );
  OR2_X1 U11255 ( .A1(n9644), .A2(n9614), .ZN(n9618) );
  INV_X1 U11256 ( .A(n11194), .ZN(n10645) );
  INV_X1 U11257 ( .A(n12798), .ZN(n11648) );
  NAND2_X1 U11258 ( .A1(n10645), .A2(n11648), .ZN(n9619) );
  NAND2_X1 U11259 ( .A1(n9984), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n9630) );
  NAND2_X1 U11260 ( .A1(n7437), .A2(n14472), .ZN(n9629) );
  INV_X1 U11261 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n9620) );
  OR2_X1 U11262 ( .A1(n7434), .A2(n9620), .ZN(n9628) );
  INV_X1 U11263 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n9621) );
  OR2_X1 U11264 ( .A1(n7436), .A2(n9621), .ZN(n9627) );
  AND4_X1 U11265 ( .A1(n9630), .A2(n9629), .A3(n9628), .A4(n9627), .ZN(n11501)
         );
  XNOR2_X1 U11266 ( .A(n9623), .B(n9622), .ZN(n10142) );
  NAND2_X1 U11267 ( .A1(n9624), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9625) );
  XNOR2_X1 U11268 ( .A(n9625), .B(P3_IR_REG_3__SCAN_IN), .ZN(n11277) );
  OAI22_X1 U11269 ( .A1(n9644), .A2(n10142), .B1(n11277), .B2(n10928), .ZN(
        n9626) );
  NAND2_X1 U11270 ( .A1(n11501), .A2(n13484), .ZN(n12805) );
  NAND4_X1 U11271 ( .A1(n9630), .A2(n9629), .A3(n9628), .A4(n9627), .ZN(n13607) );
  INV_X1 U11272 ( .A(n11630), .ZN(n12927) );
  NAND2_X1 U11273 ( .A1(n11626), .A2(n12805), .ZN(n11474) );
  NAND2_X1 U11274 ( .A1(n9984), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9636) );
  NAND2_X1 U11275 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9631) );
  NAND2_X1 U11276 ( .A1(n9663), .A2(n9631), .ZN(n11640) );
  NAND2_X1 U11277 ( .A1(n7437), .A2(n11640), .ZN(n9635) );
  INV_X1 U11278 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n11480) );
  OR2_X1 U11279 ( .A1(n7434), .A2(n11480), .ZN(n9634) );
  INV_X1 U11280 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10941) );
  XNOR2_X1 U11281 ( .A(n9638), .B(n9637), .ZN(n10144) );
  NAND2_X1 U11282 ( .A1(n9639), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9640) );
  MUX2_X1 U11283 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9640), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n9643) );
  INV_X1 U11284 ( .A(n9641), .ZN(n9642) );
  NAND2_X1 U11285 ( .A1(n9646), .A2(n11689), .ZN(n9647) );
  NAND2_X1 U11286 ( .A1(n13485), .A2(n8016), .ZN(n12806) );
  NAND2_X1 U11287 ( .A1(n11474), .A2(n7578), .ZN(n9648) );
  NAND2_X1 U11288 ( .A1(n9648), .A2(n9647), .ZN(n11938) );
  NAND2_X1 U11289 ( .A1(n10038), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n9654) );
  XNOR2_X1 U11290 ( .A(n9663), .B(P3_REG3_REG_5__SCAN_IN), .ZN(n11953) );
  NAND2_X1 U11291 ( .A1(n7437), .A2(n11953), .ZN(n9653) );
  INV_X1 U11292 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n9650) );
  OR2_X1 U11293 ( .A1(n7434), .A2(n9650), .ZN(n9652) );
  INV_X1 U11294 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10944) );
  OR2_X1 U11295 ( .A1(n7436), .A2(n10944), .ZN(n9651) );
  XNOR2_X1 U11296 ( .A(n9656), .B(n9655), .ZN(n10151) );
  NAND2_X1 U11297 ( .A1(n12759), .A2(n10151), .ZN(n9660) );
  OR2_X1 U11298 ( .A1(n9641), .A2(n14143), .ZN(n9658) );
  XNOR2_X1 U11299 ( .A(n9658), .B(n9657), .ZN(n10955) );
  NAND2_X1 U11300 ( .A1(n9768), .A2(n10955), .ZN(n9659) );
  NAND2_X1 U11301 ( .A1(n11754), .A2(n11706), .ZN(n12810) );
  INV_X1 U11302 ( .A(n11706), .ZN(n9997) );
  NAND2_X1 U11303 ( .A1(n12163), .A2(n9997), .ZN(n12809) );
  NAND2_X1 U11304 ( .A1(n11938), .A2(n12925), .ZN(n11940) );
  NAND2_X1 U11305 ( .A1(n10038), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9668) );
  NAND2_X1 U11306 ( .A1(n9954), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9667) );
  OAI21_X1 U11307 ( .B1(n9663), .B2(P3_REG3_REG_5__SCAN_IN), .A(
        P3_REG3_REG_6__SCAN_IN), .ZN(n9664) );
  NAND2_X1 U11308 ( .A1(n9664), .A2(n9675), .ZN(n12161) );
  NAND2_X1 U11309 ( .A1(n9632), .A2(n12161), .ZN(n9666) );
  NAND2_X1 U11310 ( .A1(n7435), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9665) );
  NAND2_X1 U11311 ( .A1(n12760), .A2(SI_6_), .ZN(n9674) );
  XNOR2_X1 U11312 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n9669) );
  XNOR2_X1 U11313 ( .A(n9670), .B(n9669), .ZN(n10153) );
  NAND2_X1 U11314 ( .A1(n12759), .A2(n10153), .ZN(n9673) );
  OR2_X1 U11315 ( .A1(n9686), .A2(n14143), .ZN(n9671) );
  XNOR2_X1 U11316 ( .A(n9671), .B(P3_IR_REG_6__SCAN_IN), .ZN(n11230) );
  NAND2_X1 U11317 ( .A1(n9768), .A2(n11230), .ZN(n9672) );
  XNOR2_X1 U11318 ( .A(n13605), .B(n12814), .ZN(n12931) );
  INV_X1 U11319 ( .A(n13605), .ZN(n12384) );
  NAND2_X1 U11320 ( .A1(n12384), .A2(n12164), .ZN(n12816) );
  NAND2_X1 U11321 ( .A1(n10038), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n9680) );
  NAND2_X1 U11322 ( .A1(n9675), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9676) );
  NAND2_X1 U11323 ( .A1(n9692), .A2(n9676), .ZN(n13446) );
  NAND2_X1 U11324 ( .A1(n7437), .A2(n13446), .ZN(n9679) );
  INV_X1 U11325 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n12115) );
  OR2_X1 U11326 ( .A1(n7434), .A2(n12115), .ZN(n9678) );
  INV_X1 U11327 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n12285) );
  OR2_X1 U11328 ( .A1(n7436), .A2(n12285), .ZN(n9677) );
  NAND2_X1 U11329 ( .A1(n12760), .A2(n10148), .ZN(n9691) );
  NAND2_X1 U11330 ( .A1(n9682), .A2(n9681), .ZN(n9683) );
  NAND2_X1 U11331 ( .A1(n9684), .A2(n9683), .ZN(n10147) );
  NAND2_X1 U11332 ( .A1(n12759), .A2(n10147), .ZN(n9690) );
  NAND2_X1 U11333 ( .A1(n9686), .A2(n9685), .ZN(n9700) );
  NAND2_X1 U11334 ( .A1(n9700), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9688) );
  INV_X1 U11335 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9687) );
  XNOR2_X1 U11336 ( .A(n9688), .B(n9687), .ZN(n11385) );
  NAND2_X1 U11337 ( .A1(n9768), .A2(n11385), .ZN(n9689) );
  NAND2_X1 U11338 ( .A1(n12388), .A2(n13445), .ZN(n12820) );
  INV_X1 U11339 ( .A(n13445), .ZN(n12116) );
  NAND2_X1 U11340 ( .A1(n12394), .A2(n12116), .ZN(n12819) );
  NAND2_X1 U11341 ( .A1(n12820), .A2(n12819), .ZN(n10000) );
  NAND2_X1 U11342 ( .A1(n10038), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n9697) );
  INV_X1 U11343 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11390) );
  OR2_X1 U11344 ( .A1(n7436), .A2(n11390), .ZN(n9696) );
  NAND2_X1 U11345 ( .A1(n9954), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9695) );
  NAND2_X1 U11346 ( .A1(n9692), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9693) );
  NAND2_X1 U11347 ( .A1(n9704), .A2(n9693), .ZN(n12392) );
  NAND2_X1 U11348 ( .A1(n9632), .A2(n12392), .ZN(n9694) );
  NAND4_X1 U11349 ( .A1(n9697), .A2(n9696), .A3(n9695), .A4(n9694), .ZN(n13604) );
  XNOR2_X1 U11350 ( .A(n9699), .B(n9698), .ZN(n10159) );
  NAND2_X1 U11351 ( .A1(n12760), .A2(SI_8_), .ZN(n9703) );
  NAND2_X1 U11352 ( .A1(n9715), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9701) );
  XNOR2_X1 U11353 ( .A(n9701), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11665) );
  NAND2_X1 U11354 ( .A1(n9768), .A2(n11665), .ZN(n9702) );
  OAI211_X1 U11355 ( .C1(n9644), .C2(n10159), .A(n9703), .B(n9702), .ZN(n12395) );
  XNOR2_X1 U11356 ( .A(n13604), .B(n12395), .ZN(n12932) );
  INV_X1 U11357 ( .A(n13604), .ZN(n10002) );
  NAND2_X1 U11358 ( .A1(n10002), .A2(n12395), .ZN(n12825) );
  NAND2_X1 U11359 ( .A1(n9704), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n9705) );
  NAND2_X1 U11360 ( .A1(n9722), .A2(n9705), .ZN(n12453) );
  NAND2_X1 U11361 ( .A1(n9632), .A2(n12453), .ZN(n9710) );
  NAND2_X1 U11362 ( .A1(n10038), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n9709) );
  INV_X1 U11363 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n9706) );
  OR2_X1 U11364 ( .A1(n7434), .A2(n9706), .ZN(n9708) );
  INV_X1 U11365 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11674) );
  OR2_X1 U11366 ( .A1(n7436), .A2(n11674), .ZN(n9707) );
  NAND2_X1 U11367 ( .A1(n9712), .A2(n9711), .ZN(n9713) );
  NAND2_X1 U11368 ( .A1(n9714), .A2(n9713), .ZN(n10161) );
  NAND2_X1 U11369 ( .A1(n12759), .A2(n10161), .ZN(n9721) );
  NOR2_X1 U11370 ( .A1(n9715), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n9718) );
  OR2_X1 U11371 ( .A1(n9718), .A2(n14143), .ZN(n9716) );
  INV_X1 U11372 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9717) );
  MUX2_X1 U11373 ( .A(n9716), .B(P3_IR_REG_31__SCAN_IN), .S(n9717), .Z(n9719)
         );
  NAND2_X1 U11374 ( .A1(n9718), .A2(n9717), .ZN(n9746) );
  NAND2_X1 U11375 ( .A1(n9719), .A2(n9746), .ZN(n11720) );
  NAND2_X1 U11376 ( .A1(n9768), .A2(n11720), .ZN(n9720) );
  NOR2_X1 U11377 ( .A1(n13603), .A2(n12462), .ZN(n12828) );
  NAND2_X1 U11378 ( .A1(n13603), .A2(n12462), .ZN(n12829) );
  NAND2_X1 U11379 ( .A1(n10038), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9727) );
  NAND2_X1 U11380 ( .A1(n9954), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9726) );
  NAND2_X1 U11381 ( .A1(n9722), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9723) );
  NAND2_X1 U11382 ( .A1(n9736), .A2(n9723), .ZN(n12304) );
  NAND2_X1 U11383 ( .A1(n7437), .A2(n12304), .ZN(n9725) );
  NAND2_X1 U11384 ( .A1(n7435), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n9724) );
  OAI21_X1 U11385 ( .B1(n9730), .B2(n9729), .A(n9728), .ZN(n10177) );
  NAND2_X1 U11386 ( .A1(n12759), .A2(n10177), .ZN(n9735) );
  NAND2_X1 U11387 ( .A1(n12760), .A2(n14440), .ZN(n9734) );
  NAND2_X1 U11388 ( .A1(n9746), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9732) );
  XNOR2_X1 U11389 ( .A(n9732), .B(n9731), .ZN(n11773) );
  NAND2_X1 U11390 ( .A1(n9768), .A2(n11773), .ZN(n9733) );
  XNOR2_X1 U11391 ( .A(n12832), .B(n12546), .ZN(n12934) );
  INV_X1 U11392 ( .A(n12832), .ZN(n12461) );
  NAND2_X1 U11393 ( .A1(n12461), .A2(n12546), .ZN(n12834) );
  NAND2_X1 U11394 ( .A1(n9984), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n9743) );
  NAND2_X1 U11395 ( .A1(n9736), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9737) );
  NAND2_X1 U11396 ( .A1(n9752), .A2(n9737), .ZN(n12661) );
  NAND2_X1 U11397 ( .A1(n9632), .A2(n12661), .ZN(n9742) );
  INV_X1 U11398 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n9738) );
  OR2_X1 U11399 ( .A1(n7434), .A2(n9738), .ZN(n9741) );
  INV_X1 U11400 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n9739) );
  OR2_X1 U11401 ( .A1(n7436), .A2(n9739), .ZN(n9740) );
  XNOR2_X1 U11402 ( .A(n9744), .B(n9745), .ZN(n10213) );
  NAND2_X1 U11403 ( .A1(n12759), .A2(n10213), .ZN(n9750) );
  OAI21_X1 U11404 ( .B1(n9746), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9748) );
  INV_X1 U11405 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9747) );
  XNOR2_X1 U11406 ( .A(n9748), .B(n9747), .ZN(n11904) );
  NAND2_X1 U11407 ( .A1(n9768), .A2(n11904), .ZN(n9749) );
  OAI211_X1 U11408 ( .C1(SI_11_), .C2(n7430), .A(n9750), .B(n9749), .ZN(n16581) );
  INV_X1 U11409 ( .A(n16581), .ZN(n12671) );
  NAND2_X1 U11410 ( .A1(n13971), .A2(n12671), .ZN(n12839) );
  NAND2_X1 U11411 ( .A1(n12618), .A2(n16581), .ZN(n12840) );
  NAND2_X1 U11412 ( .A1(n9984), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n9757) );
  NAND2_X1 U11413 ( .A1(n9954), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9756) );
  NAND2_X1 U11414 ( .A1(n9752), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9753) );
  NAND2_X1 U11415 ( .A1(n9781), .A2(n9753), .ZN(n13979) );
  NAND2_X1 U11416 ( .A1(n9632), .A2(n13979), .ZN(n9755) );
  NAND2_X1 U11417 ( .A1(n7435), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n9754) );
  INV_X1 U11418 ( .A(n9759), .ZN(n9760) );
  NAND2_X1 U11419 ( .A1(n8176), .A2(n9760), .ZN(n9761) );
  NAND2_X1 U11420 ( .A1(n9762), .A2(n9761), .ZN(n10230) );
  NAND2_X1 U11421 ( .A1(n12759), .A2(n10230), .ZN(n9771) );
  NAND2_X1 U11422 ( .A1(n12760), .A2(n14236), .ZN(n9770) );
  NAND2_X1 U11423 ( .A1(n9763), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9764) );
  MUX2_X1 U11424 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9764), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n9767) );
  NAND2_X1 U11425 ( .A1(n9767), .A2(n9766), .ZN(n11895) );
  NAND2_X1 U11426 ( .A1(n9768), .A2(n11895), .ZN(n9769) );
  NAND2_X1 U11427 ( .A1(n13376), .A2(n14060), .ZN(n12844) );
  INV_X1 U11428 ( .A(n14060), .ZN(n14138) );
  NAND2_X1 U11429 ( .A1(n13953), .A2(n14138), .ZN(n12843) );
  NAND2_X1 U11430 ( .A1(n13964), .A2(n13966), .ZN(n9772) );
  NAND2_X1 U11431 ( .A1(n9773), .A2(n10492), .ZN(n9774) );
  NAND2_X1 U11432 ( .A1(n9775), .A2(n9774), .ZN(n10246) );
  NAND2_X1 U11433 ( .A1(n10246), .A2(n12759), .ZN(n9780) );
  NAND2_X1 U11434 ( .A1(n9766), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9776) );
  MUX2_X1 U11435 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9776), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n9777) );
  NAND2_X1 U11436 ( .A1(n9777), .A2(n9791), .ZN(n12498) );
  INV_X1 U11437 ( .A(n12498), .ZN(n12486) );
  OAI22_X1 U11438 ( .A1(n7430), .A2(SI_13_), .B1(n12486), .B2(n10928), .ZN(
        n9778) );
  INV_X1 U11439 ( .A(n9778), .ZN(n9779) );
  NAND2_X1 U11440 ( .A1(n9954), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9786) );
  INV_X1 U11441 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13948) );
  OR2_X1 U11442 ( .A1(n7436), .A2(n13948), .ZN(n9785) );
  NAND2_X1 U11443 ( .A1(n9781), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9782) );
  NAND2_X1 U11444 ( .A1(n9796), .A2(n9782), .ZN(n13945) );
  NAND2_X1 U11445 ( .A1(n9632), .A2(n13945), .ZN(n9784) );
  NAND2_X1 U11446 ( .A1(n9984), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9783) );
  NAND4_X1 U11447 ( .A1(n9786), .A2(n9785), .A3(n9784), .A4(n9783), .ZN(n13968) );
  NAND2_X1 U11448 ( .A1(n13961), .A2(n13968), .ZN(n13930) );
  INV_X1 U11449 ( .A(n13968), .ZN(n13467) );
  NAND2_X1 U11450 ( .A1(n14055), .A2(n13467), .ZN(n9787) );
  NAND2_X1 U11451 ( .A1(n13944), .A2(n13949), .ZN(n9788) );
  NAND2_X1 U11452 ( .A1(n13961), .A2(n13467), .ZN(n12782) );
  NAND2_X1 U11453 ( .A1(n9788), .A2(n12782), .ZN(n13928) );
  XNOR2_X1 U11454 ( .A(n9789), .B(n9790), .ZN(n10383) );
  NAND2_X1 U11455 ( .A1(n10383), .A2(n12759), .ZN(n9795) );
  NAND2_X1 U11456 ( .A1(n9791), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9792) );
  XNOR2_X1 U11457 ( .A(n9792), .B(P3_IR_REG_14__SCAN_IN), .ZN(n13628) );
  OAI22_X1 U11458 ( .A1(n7430), .A2(SI_14_), .B1(n13628), .B2(n10928), .ZN(
        n9793) );
  INV_X1 U11459 ( .A(n9793), .ZN(n9794) );
  NAND2_X1 U11460 ( .A1(n10038), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9801) );
  NAND2_X1 U11461 ( .A1(n9796), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9797) );
  NAND2_X1 U11462 ( .A1(n9812), .A2(n9797), .ZN(n13937) );
  NAND2_X1 U11463 ( .A1(n9632), .A2(n13937), .ZN(n9800) );
  INV_X1 U11464 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14125) );
  OR2_X1 U11465 ( .A1(n7434), .A2(n14125), .ZN(n9799) );
  INV_X1 U11466 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13629) );
  OR2_X1 U11467 ( .A1(n7436), .A2(n13629), .ZN(n9798) );
  NAND2_X1 U11468 ( .A1(n13469), .A2(n13550), .ZN(n12785) );
  NAND2_X1 U11469 ( .A1(n14127), .A2(n13955), .ZN(n12784) );
  NAND2_X1 U11470 ( .A1(n12785), .A2(n12784), .ZN(n12848) );
  INV_X1 U11471 ( .A(n12848), .ZN(n13931) );
  NAND2_X1 U11472 ( .A1(n13928), .A2(n13931), .ZN(n9802) );
  NAND2_X1 U11473 ( .A1(n9802), .A2(n12785), .ZN(n13915) );
  NAND2_X1 U11474 ( .A1(n9804), .A2(n9803), .ZN(n9805) );
  AND2_X1 U11475 ( .A1(n9806), .A2(n9805), .ZN(n10598) );
  NAND2_X1 U11476 ( .A1(n10598), .A2(n12759), .ZN(n9811) );
  OR2_X1 U11477 ( .A1(n9807), .A2(n14143), .ZN(n9808) );
  XNOR2_X1 U11478 ( .A(n9808), .B(P3_IR_REG_15__SCAN_IN), .ZN(n13632) );
  OAI22_X1 U11479 ( .A1(n7430), .A2(n14430), .B1(n10928), .B2(n16366), .ZN(
        n9809) );
  INV_X1 U11480 ( .A(n9809), .ZN(n9810) );
  NAND2_X1 U11481 ( .A1(n9954), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9817) );
  INV_X1 U11482 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n16363) );
  OR2_X1 U11483 ( .A1(n7436), .A2(n16363), .ZN(n9816) );
  NAND2_X1 U11484 ( .A1(n9984), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n9815) );
  NAND2_X1 U11485 ( .A1(n9812), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9813) );
  NAND2_X1 U11486 ( .A1(n9832), .A2(n9813), .ZN(n13923) );
  NAND2_X1 U11487 ( .A1(n9632), .A2(n13923), .ZN(n9814) );
  NAND4_X1 U11488 ( .A1(n9817), .A2(n9816), .A3(n9815), .A4(n9814), .ZN(n13934) );
  NAND2_X1 U11489 ( .A1(n14123), .A2(n13934), .ZN(n12856) );
  INV_X1 U11490 ( .A(n13934), .ZN(n13514) );
  NAND2_X1 U11491 ( .A1(n13597), .A2(n13514), .ZN(n12855) );
  NAND2_X1 U11492 ( .A1(n12856), .A2(n12855), .ZN(n12940) );
  NAND2_X1 U11493 ( .A1(n13915), .A2(n13917), .ZN(n9818) );
  NAND2_X1 U11494 ( .A1(n9818), .A2(n12855), .ZN(n13908) );
  INV_X1 U11495 ( .A(n9819), .ZN(n9821) );
  NAND2_X1 U11496 ( .A1(n9821), .A2(n9820), .ZN(n9823) );
  AND2_X1 U11497 ( .A1(n9823), .A2(n9822), .ZN(n10656) );
  NAND2_X1 U11498 ( .A1(n10656), .A2(n12759), .ZN(n9830) );
  NAND2_X1 U11499 ( .A1(n9824), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9825) );
  MUX2_X1 U11500 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9825), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n9827) );
  NAND2_X1 U11501 ( .A1(n9827), .A2(n9840), .ZN(n13649) );
  OAI22_X1 U11502 ( .A1(n7430), .A2(n14429), .B1(n10928), .B2(n13649), .ZN(
        n9828) );
  INV_X1 U11503 ( .A(n9828), .ZN(n9829) );
  NAND2_X1 U11504 ( .A1(n10038), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n9837) );
  INV_X1 U11505 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n9831) );
  OR2_X1 U11506 ( .A1(n7436), .A2(n9831), .ZN(n9836) );
  NAND2_X1 U11507 ( .A1(n10039), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9835) );
  NAND2_X1 U11508 ( .A1(n9832), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9833) );
  NAND2_X1 U11509 ( .A1(n9846), .A2(n9833), .ZN(n13909) );
  NAND2_X1 U11510 ( .A1(n9632), .A2(n13909), .ZN(n9834) );
  NAND4_X1 U11511 ( .A1(n9837), .A2(n9836), .A3(n9835), .A4(n9834), .ZN(n13920) );
  NAND2_X1 U11512 ( .A1(n13912), .A2(n13920), .ZN(n12862) );
  NAND2_X1 U11513 ( .A1(n14039), .A2(n13594), .ZN(n12860) );
  NAND2_X1 U11514 ( .A1(n13908), .A2(n13907), .ZN(n13906) );
  NAND2_X1 U11515 ( .A1(n13906), .A2(n12860), .ZN(n13888) );
  XNOR2_X1 U11516 ( .A(n9839), .B(n9838), .ZN(n10827) );
  NAND2_X1 U11517 ( .A1(n10827), .A2(n12759), .ZN(n9845) );
  INV_X1 U11518 ( .A(SI_17_), .ZN(n10829) );
  NAND2_X1 U11519 ( .A1(n9840), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9841) );
  MUX2_X1 U11520 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9841), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n9842) );
  NAND2_X1 U11521 ( .A1(n9842), .A2(n9857), .ZN(n13668) );
  OAI22_X1 U11522 ( .A1(n7430), .A2(n10829), .B1(n10928), .B2(n13668), .ZN(
        n9843) );
  INV_X1 U11523 ( .A(n9843), .ZN(n9844) );
  NAND2_X1 U11524 ( .A1(n9984), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9851) );
  NAND2_X1 U11525 ( .A1(n9846), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9847) );
  NAND2_X1 U11526 ( .A1(n9863), .A2(n9847), .ZN(n13897) );
  NAND2_X1 U11527 ( .A1(n9632), .A2(n13897), .ZN(n9850) );
  INV_X1 U11528 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n14116) );
  OR2_X1 U11529 ( .A1(n7434), .A2(n14116), .ZN(n9849) );
  INV_X1 U11530 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13651) );
  OR2_X1 U11531 ( .A1(n7436), .A2(n13651), .ZN(n9848) );
  OR2_X1 U11532 ( .A1(n13896), .A2(n13881), .ZN(n12864) );
  NAND2_X1 U11533 ( .A1(n13896), .A2(n13881), .ZN(n12872) );
  NAND2_X1 U11534 ( .A1(n12864), .A2(n12872), .ZN(n13890) );
  NAND2_X1 U11535 ( .A1(n13888), .A2(n13887), .ZN(n9852) );
  NAND2_X1 U11536 ( .A1(n9854), .A2(n9853), .ZN(n9855) );
  NAND2_X1 U11537 ( .A1(n9856), .A2(n9855), .ZN(n10845) );
  OR2_X1 U11538 ( .A1(n10845), .A2(n9644), .ZN(n9862) );
  NAND2_X1 U11539 ( .A1(n9857), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9859) );
  INV_X1 U11540 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n9858) );
  XNOR2_X1 U11541 ( .A(n9859), .B(n9858), .ZN(n13680) );
  OAI22_X1 U11542 ( .A1(n7430), .A2(n14425), .B1(n10928), .B2(n13680), .ZN(
        n9860) );
  INV_X1 U11543 ( .A(n9860), .ZN(n9861) );
  NAND2_X1 U11544 ( .A1(n10039), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9868) );
  NAND2_X1 U11545 ( .A1(n7435), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9867) );
  NAND2_X1 U11546 ( .A1(n9863), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9864) );
  NAND2_X1 U11547 ( .A1(n9875), .A2(n9864), .ZN(n13882) );
  NAND2_X1 U11548 ( .A1(n9632), .A2(n13882), .ZN(n9866) );
  NAND2_X1 U11549 ( .A1(n9984), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9865) );
  NAND4_X1 U11550 ( .A1(n9868), .A2(n9867), .A3(n9866), .A4(n9865), .ZN(n13892) );
  NAND2_X1 U11551 ( .A1(n13884), .A2(n13892), .ZN(n12869) );
  OAI21_X1 U11552 ( .B1(n9869), .B2(n9871), .A(n9870), .ZN(n11162) );
  OR2_X1 U11553 ( .A1(n11162), .A2(n9644), .ZN(n9874) );
  OAI22_X1 U11554 ( .A1(n7430), .A2(n14424), .B1(n10928), .B2(n13694), .ZN(
        n9872) );
  INV_X1 U11555 ( .A(n9872), .ZN(n9873) );
  INV_X1 U11556 ( .A(n14027), .ZN(n13871) );
  NAND2_X1 U11557 ( .A1(n9954), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9880) );
  NAND2_X1 U11558 ( .A1(n10038), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9879) );
  NAND2_X1 U11559 ( .A1(n9875), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9876) );
  NAND2_X1 U11560 ( .A1(n9885), .A2(n9876), .ZN(n13869) );
  NAND2_X1 U11561 ( .A1(n9632), .A2(n13869), .ZN(n9878) );
  NAND2_X1 U11562 ( .A1(n7435), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n9877) );
  NAND4_X1 U11563 ( .A1(n9880), .A2(n9879), .A3(n9878), .A4(n9877), .ZN(n13856) );
  NAND2_X1 U11564 ( .A1(n13871), .A2(n13856), .ZN(n12874) );
  NAND2_X1 U11565 ( .A1(n14027), .A2(n13879), .ZN(n12871) );
  XNOR2_X1 U11566 ( .A(n9881), .B(n9882), .ZN(n11280) );
  NAND2_X1 U11567 ( .A1(n11280), .A2(n12759), .ZN(n9884) );
  NAND2_X1 U11568 ( .A1(n12760), .A2(SI_20_), .ZN(n9883) );
  NAND2_X1 U11569 ( .A1(n10038), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9892) );
  NAND2_X1 U11570 ( .A1(n9885), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9886) );
  NAND2_X1 U11571 ( .A1(n9899), .A2(n9886), .ZN(n13860) );
  NAND2_X1 U11572 ( .A1(n9632), .A2(n13860), .ZN(n9891) );
  INV_X1 U11573 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n9887) );
  OR2_X1 U11574 ( .A1(n7434), .A2(n9887), .ZN(n9890) );
  INV_X1 U11575 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n9888) );
  OR2_X1 U11576 ( .A1(n7436), .A2(n9888), .ZN(n9889) );
  NAND2_X1 U11577 ( .A1(n14023), .A2(n13867), .ZN(n12880) );
  INV_X1 U11578 ( .A(n9893), .ZN(n9894) );
  NAND2_X1 U11579 ( .A1(n7511), .A2(n9894), .ZN(n9895) );
  AND2_X1 U11580 ( .A1(n9896), .A2(n9895), .ZN(n11441) );
  NAND2_X1 U11581 ( .A1(n11441), .A2(n12759), .ZN(n9898) );
  NAND2_X1 U11582 ( .A1(n12760), .A2(SI_21_), .ZN(n9897) );
  NAND2_X1 U11583 ( .A1(n9954), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n9904) );
  NAND2_X1 U11584 ( .A1(n7435), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9903) );
  NAND2_X1 U11585 ( .A1(n9899), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9900) );
  NAND2_X1 U11586 ( .A1(n9911), .A2(n9900), .ZN(n13842) );
  NAND2_X1 U11587 ( .A1(n9632), .A2(n13842), .ZN(n9902) );
  NAND2_X1 U11588 ( .A1(n10038), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9901) );
  NAND4_X1 U11589 ( .A1(n9904), .A2(n9903), .A3(n9902), .A4(n9901), .ZN(n13855) );
  NAND2_X1 U11590 ( .A1(n14020), .A2(n13855), .ZN(n10021) );
  INV_X1 U11591 ( .A(n13855), .ZN(n13823) );
  NAND2_X1 U11592 ( .A1(n14020), .A2(n13823), .ZN(n13401) );
  XNOR2_X1 U11593 ( .A(n9906), .B(n9905), .ZN(n11496) );
  NAND2_X1 U11594 ( .A1(n11496), .A2(n12759), .ZN(n9908) );
  NAND2_X1 U11595 ( .A1(n12760), .A2(SI_22_), .ZN(n9907) );
  INV_X1 U11596 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13821) );
  NAND2_X1 U11597 ( .A1(n10038), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9910) );
  NAND2_X1 U11598 ( .A1(n9954), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n9909) );
  AND2_X1 U11599 ( .A1(n9910), .A2(n9909), .ZN(n9914) );
  NAND2_X1 U11600 ( .A1(n9911), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9912) );
  NAND2_X1 U11601 ( .A1(n9920), .A2(n9912), .ZN(n13819) );
  NAND2_X1 U11602 ( .A1(n13819), .A2(n9632), .ZN(n9913) );
  XNOR2_X1 U11603 ( .A(n14012), .B(n13833), .ZN(n13817) );
  INV_X1 U11604 ( .A(n13833), .ZN(n13806) );
  NAND2_X1 U11605 ( .A1(n14012), .A2(n13806), .ZN(n9915) );
  XNOR2_X1 U11606 ( .A(n9917), .B(n9916), .ZN(n11703) );
  NAND2_X1 U11607 ( .A1(n11703), .A2(n12759), .ZN(n9919) );
  NAND2_X1 U11608 ( .A1(n12760), .A2(SI_23_), .ZN(n9918) );
  NAND2_X1 U11609 ( .A1(n9920), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9921) );
  NAND2_X1 U11610 ( .A1(n9928), .A2(n9921), .ZN(n13812) );
  NAND2_X1 U11611 ( .A1(n13812), .A2(n9632), .ZN(n9924) );
  AOI22_X1 U11612 ( .A1(n9984), .A2(P3_REG1_REG_23__SCAN_IN), .B1(n10039), 
        .B2(P3_REG0_REG_23__SCAN_IN), .ZN(n9923) );
  NAND2_X1 U11613 ( .A1(n7435), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9922) );
  XNOR2_X1 U11614 ( .A(n9925), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n12257) );
  NAND2_X1 U11615 ( .A1(n12257), .A2(n12759), .ZN(n9927) );
  NAND2_X1 U11616 ( .A1(n12760), .A2(SI_24_), .ZN(n9926) );
  INV_X1 U11617 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n13798) );
  NAND2_X1 U11618 ( .A1(n9928), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9929) );
  NAND2_X1 U11619 ( .A1(n9939), .A2(n9929), .ZN(n13800) );
  NAND2_X1 U11620 ( .A1(n13800), .A2(n9632), .ZN(n9931) );
  AOI22_X1 U11621 ( .A1(n9984), .A2(P3_REG1_REG_24__SCAN_IN), .B1(n10039), 
        .B2(P3_REG0_REG_24__SCAN_IN), .ZN(n9930) );
  OAI211_X1 U11622 ( .C1(n7436), .C2(n13798), .A(n9931), .B(n9930), .ZN(n13602) );
  NAND2_X1 U11623 ( .A1(n13801), .A2(n13807), .ZN(n12780) );
  NAND2_X1 U11624 ( .A1(n9934), .A2(n9933), .ZN(n9936) );
  NAND2_X1 U11625 ( .A1(n9936), .A2(n9935), .ZN(n12350) );
  NAND2_X1 U11626 ( .A1(n12760), .A2(SI_25_), .ZN(n9937) );
  NAND2_X1 U11627 ( .A1(n9939), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9940) );
  NAND2_X1 U11628 ( .A1(n9952), .A2(n9940), .ZN(n13784) );
  NAND2_X1 U11629 ( .A1(n13784), .A2(n9632), .ZN(n9945) );
  INV_X1 U11630 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n13785) );
  NAND2_X1 U11631 ( .A1(n9954), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n9942) );
  NAND2_X1 U11632 ( .A1(n9984), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9941) );
  OAI211_X1 U11633 ( .C1(n7436), .C2(n13785), .A(n9942), .B(n9941), .ZN(n9943)
         );
  INV_X1 U11634 ( .A(n9943), .ZN(n9944) );
  NAND2_X1 U11635 ( .A1(n14001), .A2(n13531), .ZN(n12768) );
  NAND2_X1 U11636 ( .A1(n13776), .A2(n12768), .ZN(n9946) );
  NAND2_X1 U11637 ( .A1(n13507), .A2(n13795), .ZN(n10029) );
  NAND2_X1 U11638 ( .A1(n9946), .A2(n10029), .ZN(n13763) );
  OR2_X1 U11639 ( .A1(n9948), .A2(n9947), .ZN(n9950) );
  NAND2_X1 U11640 ( .A1(n12760), .A2(SI_26_), .ZN(n9951) );
  NAND2_X1 U11641 ( .A1(n9952), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9953) );
  NAND2_X1 U11642 ( .A1(n9967), .A2(n9953), .ZN(n13773) );
  NAND2_X1 U11643 ( .A1(n13773), .A2(n9632), .ZN(n9959) );
  INV_X1 U11644 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n13772) );
  NAND2_X1 U11645 ( .A1(n10038), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9956) );
  NAND2_X1 U11646 ( .A1(n9954), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9955) );
  OAI211_X1 U11647 ( .C1(n13772), .C2(n7436), .A(n9956), .B(n9955), .ZN(n9957)
         );
  INV_X1 U11648 ( .A(n9957), .ZN(n9958) );
  NAND2_X1 U11649 ( .A1(n13996), .A2(n13779), .ZN(n12769) );
  NAND2_X1 U11650 ( .A1(n13763), .A2(n12769), .ZN(n9960) );
  NAND2_X1 U11651 ( .A1(n9960), .A2(n12771), .ZN(n13746) );
  NAND2_X1 U11652 ( .A1(n12760), .A2(SI_27_), .ZN(n9965) );
  NAND2_X1 U11653 ( .A1(n9967), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9968) );
  NAND2_X1 U11654 ( .A1(n9982), .A2(n9968), .ZN(n13758) );
  NAND2_X1 U11655 ( .A1(n13758), .A2(n9632), .ZN(n9974) );
  INV_X1 U11656 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n9971) );
  NAND2_X1 U11657 ( .A1(n10038), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9970) );
  NAND2_X1 U11658 ( .A1(n9954), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9969) );
  OAI211_X1 U11659 ( .C1(n9971), .C2(n7436), .A(n9970), .B(n9969), .ZN(n9972)
         );
  INV_X1 U11660 ( .A(n9972), .ZN(n9973) );
  NAND2_X2 U11661 ( .A1(n9974), .A2(n9973), .ZN(n13768) );
  XNOR2_X2 U11662 ( .A(n13759), .B(n13768), .ZN(n13750) );
  NAND2_X1 U11663 ( .A1(n13746), .A2(n13750), .ZN(n9975) );
  NAND2_X1 U11664 ( .A1(n14076), .A2(n13768), .ZN(n12772) );
  NAND2_X1 U11665 ( .A1(n9975), .A2(n12772), .ZN(n13742) );
  OR2_X1 U11666 ( .A1(n9977), .A2(n9976), .ZN(n9978) );
  NAND2_X1 U11667 ( .A1(n9979), .A2(n9978), .ZN(n12733) );
  NAND2_X1 U11668 ( .A1(n12760), .A2(SI_28_), .ZN(n9980) );
  NAND2_X1 U11669 ( .A1(n9982), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9983) );
  NAND2_X1 U11670 ( .A1(n13718), .A2(n9983), .ZN(n13431) );
  INV_X1 U11671 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n13738) );
  NAND2_X1 U11672 ( .A1(n9984), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9986) );
  NAND2_X1 U11673 ( .A1(n10039), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9985) );
  OAI211_X1 U11674 ( .C1(n13738), .C2(n7436), .A(n9986), .B(n9985), .ZN(n9987)
         );
  AOI21_X2 U11675 ( .B1(n13431), .B2(n9632), .A(n9987), .ZN(n13754) );
  OR2_X2 U11676 ( .A1(n13741), .A2(n13754), .ZN(n12908) );
  NAND2_X1 U11677 ( .A1(n13741), .A2(n13754), .ZN(n9988) );
  NAND2_X2 U11678 ( .A1(n12908), .A2(n9988), .ZN(n13743) );
  INV_X1 U11679 ( .A(n13743), .ZN(n12899) );
  INV_X1 U11680 ( .A(n12908), .ZN(n9989) );
  INV_X1 U11681 ( .A(n13741), .ZN(n14074) );
  NAND2_X1 U11682 ( .A1(n10636), .A2(n11032), .ZN(n11031) );
  NAND2_X1 U11683 ( .A1(n12922), .A2(n11031), .ZN(n11530) );
  NAND2_X1 U11684 ( .A1(n11654), .A2(n11529), .ZN(n9991) );
  NAND2_X1 U11685 ( .A1(n11530), .A2(n9991), .ZN(n11653) );
  NAND2_X1 U11686 ( .A1(n11653), .A2(n12930), .ZN(n11652) );
  NAND2_X1 U11687 ( .A1(n10645), .A2(n12798), .ZN(n11629) );
  AND2_X1 U11688 ( .A1(n11630), .A2(n11629), .ZN(n9992) );
  NAND2_X1 U11689 ( .A1(n13607), .A2(n13484), .ZN(n11475) );
  NAND2_X1 U11690 ( .A1(n13485), .A2(n11689), .ZN(n9994) );
  AND2_X1 U11691 ( .A1(n11475), .A2(n9994), .ZN(n11941) );
  INV_X1 U11692 ( .A(n12925), .ZN(n9993) );
  NAND2_X1 U11693 ( .A1(n11754), .A2(n9997), .ZN(n11750) );
  AND2_X1 U11694 ( .A1(n12931), .A2(n11750), .ZN(n9998) );
  NAND2_X1 U11695 ( .A1(n11749), .A2(n9998), .ZN(n11752) );
  NAND2_X1 U11696 ( .A1(n13605), .A2(n12164), .ZN(n9999) );
  NAND2_X1 U11697 ( .A1(n11752), .A2(n9999), .ZN(n12107) );
  NAND2_X1 U11698 ( .A1(n12394), .A2(n13445), .ZN(n10001) );
  INV_X1 U11699 ( .A(n12395), .ZN(n12823) );
  NAND2_X1 U11700 ( .A1(n10002), .A2(n12823), .ZN(n10003) );
  NAND2_X1 U11701 ( .A1(n12291), .A2(n12462), .ZN(n10004) );
  NAND2_X1 U11702 ( .A1(n10005), .A2(n10004), .ZN(n12300) );
  NAND2_X1 U11703 ( .A1(n12832), .A2(n12546), .ZN(n10007) );
  NAND2_X1 U11704 ( .A1(n13971), .A2(n16581), .ZN(n10008) );
  NAND2_X1 U11705 ( .A1(n12618), .A2(n12671), .ZN(n10009) );
  INV_X1 U11706 ( .A(n13965), .ZN(n10010) );
  NAND2_X1 U11707 ( .A1(n13376), .A2(n14138), .ZN(n10011) );
  NAND2_X1 U11708 ( .A1(n13929), .A2(n13930), .ZN(n10013) );
  NAND2_X1 U11709 ( .A1(n13469), .A2(n13955), .ZN(n13916) );
  NAND2_X1 U11710 ( .A1(n13933), .A2(n13916), .ZN(n10014) );
  NAND2_X1 U11711 ( .A1(n13597), .A2(n13934), .ZN(n10015) );
  NAND2_X1 U11712 ( .A1(n13912), .A2(n13594), .ZN(n13891) );
  AND2_X1 U11713 ( .A1(n13890), .A2(n13891), .ZN(n10017) );
  NAND2_X1 U11714 ( .A1(n13902), .A2(n10017), .ZN(n13889) );
  NAND2_X1 U11715 ( .A1(n13896), .A2(n13904), .ZN(n10018) );
  NOR2_X1 U11716 ( .A1(n14027), .A2(n13856), .ZN(n10020) );
  AND2_X1 U11717 ( .A1(n13852), .A2(n13402), .ZN(n10026) );
  INV_X1 U11718 ( .A(n13402), .ZN(n10025) );
  NAND2_X1 U11719 ( .A1(n14023), .A2(n13834), .ZN(n13830) );
  INV_X1 U11720 ( .A(n13830), .ZN(n10023) );
  INV_X1 U11721 ( .A(n10021), .ZN(n10022) );
  NOR2_X1 U11722 ( .A1(n10023), .A2(n10022), .ZN(n10024) );
  NAND2_X1 U11723 ( .A1(n14012), .A2(n13833), .ZN(n10027) );
  AND2_X1 U11724 ( .A1(n13801), .A2(n13602), .ZN(n10028) );
  NAND2_X1 U11725 ( .A1(n14001), .A2(n13795), .ZN(n10030) );
  NAND2_X1 U11726 ( .A1(n14081), .A2(n13779), .ZN(n10031) );
  NAND2_X1 U11727 ( .A1(n13996), .A2(n13421), .ZN(n10032) );
  NAND2_X1 U11728 ( .A1(n14076), .A2(n13733), .ZN(n10034) );
  AND2_X2 U11729 ( .A1(n13748), .A2(n10034), .ZN(n13732) );
  OAI21_X1 U11730 ( .B1(n13754), .B2(n14074), .A(n13731), .ZN(n10035) );
  XNOR2_X1 U11731 ( .A(n10035), .B(n12948), .ZN(n10049) );
  INV_X1 U11732 ( .A(n11281), .ZN(n10095) );
  NAND2_X1 U11733 ( .A1(n12789), .A2(n10095), .ZN(n12763) );
  INV_X1 U11734 ( .A(n12732), .ZN(n12960) );
  NAND2_X1 U11735 ( .A1(n12960), .A2(n13697), .ZN(n10930) );
  NAND2_X1 U11736 ( .A1(n10930), .A2(n10928), .ZN(n11037) );
  NAND2_X1 U11737 ( .A1(n12960), .A2(P3_B_REG_SCAN_IN), .ZN(n10037) );
  NAND2_X1 U11738 ( .A1(n13967), .A2(n10037), .ZN(n13716) );
  INV_X1 U11739 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n10042) );
  NAND2_X1 U11740 ( .A1(n10038), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n10041) );
  NAND2_X1 U11741 ( .A1(n10039), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n10040) );
  OAI211_X1 U11742 ( .C1(n10042), .C2(n7436), .A(n10041), .B(n10040), .ZN(
        n10043) );
  INV_X1 U11743 ( .A(n10043), .ZN(n10044) );
  NOR2_X1 U11744 ( .A1(n13716), .A2(n12913), .ZN(n10047) );
  INV_X1 U11745 ( .A(n11037), .ZN(n10045) );
  NAND2_X1 U11746 ( .A1(n10050), .A2(n12901), .ZN(n11516) );
  NAND2_X1 U11747 ( .A1(n10094), .A2(n12910), .ZN(n11513) );
  NAND2_X1 U11748 ( .A1(n11516), .A2(n11513), .ZN(n10062) );
  NAND2_X1 U11749 ( .A1(n10051), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10052) );
  MUX2_X1 U11750 ( .A(P3_IR_REG_31__SCAN_IN), .B(n10052), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n10054) );
  NAND2_X1 U11751 ( .A1(n10054), .A2(n10053), .ZN(n12260) );
  XNOR2_X1 U11752 ( .A(n12260), .B(P3_B_REG_SCAN_IN), .ZN(n10057) );
  NAND2_X1 U11753 ( .A1(n10053), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10055) );
  MUX2_X1 U11754 ( .A(P3_IR_REG_31__SCAN_IN), .B(n10055), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n10056) );
  NAND2_X1 U11755 ( .A1(n10056), .A2(n7468), .ZN(n12348) );
  NAND2_X1 U11756 ( .A1(n10057), .A2(n12348), .ZN(n10059) );
  NAND2_X1 U11757 ( .A1(n7468), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10058) );
  INV_X1 U11758 ( .A(n10079), .ZN(n12483) );
  NAND2_X1 U11759 ( .A1(n12483), .A2(n12348), .ZN(n10060) );
  NAND2_X1 U11760 ( .A1(n10062), .A2(n14141), .ZN(n10086) );
  NAND2_X1 U11761 ( .A1(n12483), .A2(n12260), .ZN(n11026) );
  NAND2_X1 U11762 ( .A1(n11028), .A2(n11026), .ZN(n10099) );
  XNOR2_X1 U11763 ( .A(n14141), .B(n10099), .ZN(n10081) );
  NOR2_X1 U11764 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n10066) );
  NOR4_X1 U11765 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n10065) );
  NOR4_X1 U11766 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n10064) );
  NOR4_X1 U11767 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n10063) );
  NAND4_X1 U11768 ( .A1(n10066), .A2(n10065), .A3(n10064), .A4(n10063), .ZN(
        n10072) );
  NOR4_X1 U11769 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n10070) );
  NOR4_X1 U11770 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n10069) );
  NOR4_X1 U11771 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n10068) );
  NOR4_X1 U11772 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n10067) );
  NAND4_X1 U11773 ( .A1(n10070), .A2(n10069), .A3(n10068), .A4(n10067), .ZN(
        n10071) );
  NOR2_X1 U11774 ( .A1(n10072), .A2(n10071), .ZN(n10073) );
  NOR2_X1 U11775 ( .A1(n10237), .A2(n10073), .ZN(n10098) );
  INV_X1 U11776 ( .A(n12348), .ZN(n10078) );
  INV_X1 U11777 ( .A(n12260), .ZN(n10077) );
  NAND3_X1 U11778 ( .A1(n10079), .A2(n10078), .A3(n10077), .ZN(n10737) );
  NOR2_X1 U11779 ( .A1(n10098), .A2(n10929), .ZN(n10080) );
  NAND2_X1 U11780 ( .A1(n10082), .A2(n11442), .ZN(n10083) );
  INV_X1 U11781 ( .A(n14141), .ZN(n11514) );
  OAI211_X1 U11782 ( .C1(n12963), .C2(n10084), .A(n10083), .B(n11514), .ZN(
        n10085) );
  INV_X1 U11783 ( .A(n10088), .ZN(n13727) );
  NAND2_X1 U11784 ( .A1(n10091), .A2(n10090), .ZN(P3_U3488) );
  INV_X1 U11785 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n10105) );
  INV_X1 U11786 ( .A(n10099), .ZN(n10093) );
  INV_X1 U11787 ( .A(n10098), .ZN(n10092) );
  AND3_X1 U11788 ( .A1(n10093), .A2(n10092), .A3(n14141), .ZN(n10743) );
  OR2_X1 U11789 ( .A1(n10094), .A2(n12901), .ZN(n11165) );
  NAND2_X1 U11790 ( .A1(n11442), .A2(n10095), .ZN(n12953) );
  OR2_X1 U11791 ( .A1(n10096), .A2(n12953), .ZN(n10738) );
  NAND2_X1 U11792 ( .A1(n11165), .A2(n10738), .ZN(n10097) );
  NAND2_X1 U11793 ( .A1(n10743), .A2(n10097), .ZN(n10102) );
  NOR2_X1 U11794 ( .A1(n14141), .A2(n10098), .ZN(n10100) );
  NAND2_X1 U11795 ( .A1(n10100), .A2(n10099), .ZN(n10746) );
  INV_X1 U11796 ( .A(n10728), .ZN(n10742) );
  OR2_X1 U11797 ( .A1(n10746), .A2(n10742), .ZN(n10101) );
  NAND2_X1 U11798 ( .A1(n10102), .A2(n10101), .ZN(n10103) );
  INV_X1 U11799 ( .A(n10929), .ZN(n10732) );
  NAND2_X1 U11800 ( .A1(n10088), .A2(n10106), .ZN(n10107) );
  NAND2_X1 U11801 ( .A1(n10108), .A2(n10107), .ZN(P3_U3456) );
  NOR2_X1 U11802 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), 
        .ZN(n10111) );
  NOR2_X2 U11803 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n10170) );
  NOR2_X1 U11804 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n10114) );
  INV_X1 U11805 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n10118) );
  NAND2_X1 U11806 ( .A1(n10216), .A2(n10118), .ZN(n10119) );
  NAND2_X1 U11807 ( .A1(n10215), .A2(n10214), .ZN(n10120) );
  NAND2_X1 U11808 ( .A1(n10120), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10122) );
  INV_X1 U11809 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10121) );
  NOR2_X1 U11810 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n10127) );
  NOR2_X1 U11811 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n10126) );
  NOR2_X1 U11812 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), 
        .ZN(n10125) );
  NOR2_X1 U11813 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n10124) );
  NAND2_X1 U11814 ( .A1(n10134), .A2(n10130), .ZN(n10135) );
  NAND2_X1 U11815 ( .A1(n10135), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10128) );
  MUX2_X1 U11816 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10128), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n10133) );
  NAND2_X1 U11817 ( .A1(n10136), .A2(n10135), .ZN(n15991) );
  NAND2_X1 U11818 ( .A1(n10132), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10138) );
  XNOR2_X1 U11819 ( .A(n10138), .B(n10137), .ZN(n15995) );
  NOR2_X1 U11820 ( .A1(n15991), .A2(n15995), .ZN(n10139) );
  NOR2_X1 U11821 ( .A1(n10410), .A2(P1_U3086), .ZN(n10140) );
  AND2_X2 U11822 ( .A1(n10411), .A2(n10140), .ZN(P1_U4016) );
  INV_X1 U11823 ( .A(n10737), .ZN(n10141) );
  INV_X2 U11824 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  OR3_X2 U11825 ( .A1(n10273), .A2(n10272), .A3(P2_U3088), .ZN(n14736) );
  INV_X1 U11826 ( .A(n14736), .ZN(P2_U3947) );
  AND2_X1 U11827 ( .A1(n10165), .A2(P3_U3151), .ZN(n11702) );
  AND2_X1 U11828 ( .A1(n10468), .A2(P3_U3151), .ZN(n14146) );
  AOI222_X1 U11829 ( .A1(n10142), .A2(n11702), .B1(n11277), .B2(
        P3_STATE_REG_SCAN_IN), .C1(n14146), .C2(SI_3_), .ZN(n10143) );
  INV_X1 U11830 ( .A(n10143), .ZN(P3_U3292) );
  AOI222_X1 U11831 ( .A1(n10144), .A2(n11702), .B1(n10953), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_4_), .C2(n14146), .ZN(n10145) );
  INV_X1 U11832 ( .A(n10145), .ZN(P3_U3291) );
  AND2_X1 U11833 ( .A1(n10165), .A2(P2_U3088), .ZN(n11163) );
  INV_X2 U11834 ( .A(n11163), .ZN(n15133) );
  NAND2_X1 U11835 ( .A1(n10468), .A2(P2_U3088), .ZN(n15123) );
  OAI222_X1 U11836 ( .A1(n15133), .A2(n10146), .B1(n16045), .B2(P2_U3088), 
        .C1(n15123), .C2(n10467), .ZN(P2_U3326) );
  INV_X2 U11837 ( .A(n14146), .ZN(n14150) );
  OAI222_X1 U11838 ( .A1(P3_U3151), .A2(n11385), .B1(n14150), .B2(n10148), 
        .C1(n14154), .C2(n10147), .ZN(P3_U3288) );
  OAI222_X1 U11839 ( .A1(P3_U3151), .A2(n7619), .B1(n14150), .B2(n10150), .C1(
        n14154), .C2(n10149), .ZN(P3_U3293) );
  OAI222_X1 U11840 ( .A1(P3_U3151), .A2(n10955), .B1(n14150), .B2(n10152), 
        .C1(n14154), .C2(n10151), .ZN(P3_U3290) );
  INV_X1 U11841 ( .A(n11230), .ZN(n11226) );
  INV_X2 U11842 ( .A(n11702), .ZN(n14154) );
  INV_X1 U11843 ( .A(n10153), .ZN(n10155) );
  INV_X1 U11844 ( .A(SI_6_), .ZN(n10154) );
  OAI222_X1 U11845 ( .A1(P3_U3151), .A2(n11226), .B1(n14154), .B2(n10155), 
        .C1(n10154), .C2(n14150), .ZN(P3_U3289) );
  INV_X1 U11846 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n11152) );
  INV_X1 U11847 ( .A(n10156), .ZN(n10157) );
  OAI222_X1 U11848 ( .A1(P3_U3151), .A2(n11152), .B1(n14154), .B2(n10157), 
        .C1(n10339), .C2(n14150), .ZN(P3_U3295) );
  INV_X1 U11849 ( .A(SI_8_), .ZN(n10158) );
  INV_X1 U11850 ( .A(n11665), .ZN(n11392) );
  OAI222_X1 U11851 ( .A1(n14154), .A2(n10159), .B1(n14150), .B2(n10158), .C1(
        P3_U3151), .C2(n11392), .ZN(P3_U3287) );
  INV_X1 U11852 ( .A(n10754), .ZN(n10187) );
  OAI222_X1 U11853 ( .A1(n15133), .A2(n10160), .B1(n15123), .B2(n10187), .C1(
        P2_U3088), .C2(n10287), .ZN(P2_U3323) );
  INV_X1 U11854 ( .A(SI_9_), .ZN(n10162) );
  OAI222_X1 U11855 ( .A1(P3_U3151), .A2(n11720), .B1(n14150), .B2(n10162), 
        .C1(n14154), .C2(n10161), .ZN(P3_U3286) );
  INV_X1 U11856 ( .A(n14745), .ZN(n10163) );
  INV_X1 U11857 ( .A(n10516), .ZN(n10168) );
  OAI222_X1 U11858 ( .A1(n15133), .A2(n10164), .B1(n10163), .B2(P2_U3088), 
        .C1(n15123), .C2(n10168), .ZN(P2_U3324) );
  NAND2_X1 U11859 ( .A1(n10468), .A2(P1_U3086), .ZN(n15992) );
  INV_X1 U11860 ( .A(n15992), .ZN(n15971) );
  INV_X1 U11861 ( .A(n15971), .ZN(n15987) );
  AND2_X1 U11862 ( .A1(n10165), .A2(P1_U3086), .ZN(n12468) );
  INV_X2 U11863 ( .A(n12468), .ZN(n15990) );
  INV_X1 U11864 ( .A(n10166), .ZN(n10200) );
  NAND2_X1 U11865 ( .A1(n10200), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10167) );
  XNOR2_X1 U11866 ( .A(n10167), .B(P1_IR_REG_3__SCAN_IN), .ZN(n15412) );
  OAI222_X1 U11867 ( .A1(n15987), .A2(n7671), .B1(n15990), .B2(n10168), .C1(
        P1_U3086), .C2(n7670), .ZN(P1_U3352) );
  INV_X1 U11868 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10469) );
  NAND2_X1 U11869 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n10169) );
  INV_X1 U11870 ( .A(n10170), .ZN(n10198) );
  NAND2_X1 U11871 ( .A1(n10171), .A2(n10198), .ZN(n10471) );
  OAI222_X1 U11872 ( .A1(n15987), .A2(n10469), .B1(n15990), .B2(n10467), .C1(
        P1_U3086), .C2(n10471), .ZN(P1_U3354) );
  INV_X1 U11873 ( .A(n15123), .ZN(n12470) );
  INV_X1 U11874 ( .A(n10494), .ZN(n10202) );
  INV_X1 U11875 ( .A(n10282), .ZN(n16057) );
  OAI222_X1 U11876 ( .A1(n15131), .A2(n10202), .B1(n16057), .B2(P2_U3088), 
        .C1(n10172), .C2(n15133), .ZN(P2_U3325) );
  INV_X1 U11877 ( .A(n14769), .ZN(n10174) );
  OAI222_X1 U11878 ( .A1(n15131), .A2(n10892), .B1(n10174), .B2(P2_U3088), 
        .C1(n10173), .C2(n15133), .ZN(P2_U3321) );
  INV_X1 U11879 ( .A(n10784), .ZN(n10196) );
  INV_X1 U11880 ( .A(n14756), .ZN(n10176) );
  OAI222_X1 U11881 ( .A1(n15131), .A2(n10196), .B1(n10176), .B2(P2_U3088), 
        .C1(n10175), .C2(n15133), .ZN(P2_U3322) );
  OAI222_X1 U11882 ( .A1(P3_U3151), .A2(n11773), .B1(n14150), .B2(n14440), 
        .C1(n14154), .C2(n10177), .ZN(P3_U3285) );
  AOI22_X1 U11883 ( .A1(n14797), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n11163), .ZN(n10178) );
  OAI21_X1 U11884 ( .B1(n11290), .B2(n15131), .A(n10178), .ZN(P2_U3319) );
  INV_X1 U11885 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10184) );
  NAND2_X1 U11886 ( .A1(n10411), .A2(n10179), .ZN(n10424) );
  NAND2_X1 U11887 ( .A1(n15991), .A2(P1_B_REG_SCAN_IN), .ZN(n10180) );
  MUX2_X1 U11888 ( .A(P1_B_REG_SCAN_IN), .B(n10180), .S(n15995), .Z(n10181) );
  INV_X1 U11889 ( .A(n10181), .ZN(n10182) );
  OR2_X1 U11890 ( .A1(n10424), .A2(n10401), .ZN(n16000) );
  INV_X1 U11891 ( .A(n10411), .ZN(n10223) );
  INV_X1 U11892 ( .A(n15995), .ZN(n10390) );
  NOR4_X1 U11893 ( .A1(n10223), .A2(n10391), .A3(n10390), .A4(P1_U3086), .ZN(
        n10183) );
  AOI21_X1 U11894 ( .B1(n10184), .B2(n16000), .A(n10183), .ZN(P1_U3445) );
  NAND2_X1 U11895 ( .A1(n10189), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10185) );
  XNOR2_X1 U11896 ( .A(n10185), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10755) );
  INV_X1 U11897 ( .A(n10755), .ZN(n10188) );
  OAI222_X1 U11898 ( .A1(n10188), .A2(P1_U3086), .B1(n15990), .B2(n10187), 
        .C1(n10186), .C2(n15987), .ZN(P1_U3351) );
  INV_X1 U11899 ( .A(n10189), .ZN(n10190) );
  NAND2_X1 U11900 ( .A1(n10190), .A2(n14583), .ZN(n10193) );
  NAND2_X1 U11901 ( .A1(n10203), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10191) );
  XNOR2_X1 U11902 ( .A(n10191), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10893) );
  INV_X1 U11903 ( .A(n10893), .ZN(n10444) );
  OAI222_X1 U11904 ( .A1(P1_U3086), .A2(n10444), .B1(n15990), .B2(n10892), 
        .C1(n10192), .C2(n15987), .ZN(P1_U3349) );
  NAND2_X1 U11905 ( .A1(n10193), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10194) );
  XNOR2_X1 U11906 ( .A(n10194), .B(P1_IR_REG_5__SCAN_IN), .ZN(n15431) );
  INV_X1 U11907 ( .A(n15431), .ZN(n10197) );
  OAI222_X1 U11908 ( .A1(P1_U3086), .A2(n10197), .B1(n15990), .B2(n10196), 
        .C1(n10195), .C2(n15987), .ZN(P1_U3350) );
  NAND2_X1 U11909 ( .A1(n10198), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10199) );
  MUX2_X1 U11910 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10199), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n10201) );
  NAND2_X1 U11911 ( .A1(n10201), .A2(n10200), .ZN(n15404) );
  OAI222_X1 U11912 ( .A1(P1_U3086), .A2(n15404), .B1(n15990), .B2(n10202), 
        .C1(n10493), .C2(n15987), .ZN(P1_U3353) );
  NAND2_X1 U11913 ( .A1(n10250), .A2(n14587), .ZN(n10210) );
  NAND2_X1 U11914 ( .A1(n10210), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10204) );
  XNOR2_X1 U11915 ( .A(n10204), .B(P1_IR_REG_7__SCAN_IN), .ZN(n15443) );
  INV_X1 U11916 ( .A(n15443), .ZN(n10206) );
  INV_X1 U11917 ( .A(n11060), .ZN(n10208) );
  OAI222_X1 U11918 ( .A1(n10206), .A2(P1_U3086), .B1(n15990), .B2(n10208), 
        .C1(n10205), .C2(n15992), .ZN(P1_U3348) );
  INV_X1 U11919 ( .A(n14783), .ZN(n10207) );
  OAI222_X1 U11920 ( .A1(n15133), .A2(n10209), .B1(n15123), .B2(n10208), .C1(
        P2_U3088), .C2(n10207), .ZN(P2_U3320) );
  NAND2_X1 U11921 ( .A1(n10225), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10211) );
  XNOR2_X1 U11922 ( .A(n10211), .B(P1_IR_REG_8__SCAN_IN), .ZN(n15462) );
  INV_X1 U11923 ( .A(n15462), .ZN(n10544) );
  INV_X1 U11924 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10212) );
  OAI222_X1 U11925 ( .A1(P1_U3086), .A2(n10544), .B1(n15990), .B2(n11290), 
        .C1(n10212), .C2(n15987), .ZN(P1_U3347) );
  OAI222_X1 U11926 ( .A1(P3_U3151), .A2(n11904), .B1(n14150), .B2(n14235), 
        .C1(n14154), .C2(n10213), .ZN(P3_U3284) );
  INV_X1 U11927 ( .A(n12995), .ZN(n10222) );
  XNOR2_X2 U11928 ( .A(n10221), .B(n10220), .ZN(n15982) );
  AOI21_X1 U11929 ( .B1(n10222), .B2(n10411), .A(n13154), .ZN(n10319) );
  INV_X1 U11930 ( .A(n10319), .ZN(n10224) );
  NAND2_X1 U11931 ( .A1(n10223), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13369) );
  NAND2_X1 U11932 ( .A1(n13369), .A2(n10424), .ZN(n10318) );
  AND2_X1 U11933 ( .A1(n10224), .A2(n10318), .ZN(n16162) );
  NOR2_X1 U11934 ( .A1(n16162), .A2(P1_U4016), .ZN(P1_U3085) );
  NAND2_X1 U11935 ( .A1(n10232), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10226) );
  XNOR2_X1 U11936 ( .A(n10226), .B(P1_IR_REG_9__SCAN_IN), .ZN(n15478) );
  INV_X1 U11937 ( .A(n15478), .ZN(n10545) );
  INV_X1 U11938 ( .A(n11416), .ZN(n10228) );
  OAI222_X1 U11939 ( .A1(n10545), .A2(P1_U3086), .B1(n15990), .B2(n10228), 
        .C1(n10227), .C2(n15992), .ZN(P1_U3346) );
  INV_X1 U11940 ( .A(n16151), .ZN(n10304) );
  OAI222_X1 U11941 ( .A1(n15133), .A2(n10229), .B1(n15123), .B2(n10228), .C1(
        P2_U3088), .C2(n10304), .ZN(P2_U3318) );
  OAI222_X1 U11942 ( .A1(P3_U3151), .A2(n11895), .B1(n14150), .B2(n14236), 
        .C1(n14154), .C2(n10230), .ZN(P3_U3283) );
  INV_X1 U11943 ( .A(n11585), .ZN(n10236) );
  INV_X1 U11944 ( .A(n10372), .ZN(n10314) );
  OAI222_X1 U11945 ( .A1(n15133), .A2(n10231), .B1(n15123), .B2(n10236), .C1(
        P2_U3088), .C2(n10314), .ZN(P2_U3317) );
  INV_X1 U11946 ( .A(n10232), .ZN(n10233) );
  INV_X1 U11947 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n14592) );
  NAND2_X1 U11948 ( .A1(n10233), .A2(n14592), .ZN(n10242) );
  NAND2_X1 U11949 ( .A1(n10242), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10234) );
  XNOR2_X1 U11950 ( .A(n10234), .B(P1_IR_REG_10__SCAN_IN), .ZN(n15492) );
  INV_X1 U11951 ( .A(n15492), .ZN(n15489) );
  OAI222_X1 U11952 ( .A1(n15489), .A2(P1_U3086), .B1(n15990), .B2(n10236), 
        .C1(n10235), .C2(n15987), .ZN(P1_U3345) );
  INV_X1 U11953 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n10239) );
  INV_X1 U11954 ( .A(n11026), .ZN(n10238) );
  AOI22_X1 U11955 ( .A1(n10241), .A2(n10239), .B1(n14140), .B2(n10238), .ZN(
        P3_U3376) );
  INV_X1 U11956 ( .A(n11862), .ZN(n10245) );
  AOI22_X1 U11957 ( .A1(n10576), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n11163), .ZN(n10240) );
  OAI21_X1 U11958 ( .B1(n10245), .B2(n15131), .A(n10240), .ZN(P2_U3316) );
  AND2_X1 U11959 ( .A1(n10241), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U11960 ( .A1(n10241), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U11961 ( .A1(n10241), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U11962 ( .A1(n10241), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U11963 ( .A1(n10241), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U11964 ( .A1(n10241), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U11965 ( .A1(n10241), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U11966 ( .A1(n10241), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U11967 ( .A1(n10241), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U11968 ( .A1(n10241), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U11969 ( .A1(n10241), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U11970 ( .A1(n10241), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U11971 ( .A1(n10241), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U11972 ( .A1(n10241), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U11973 ( .A1(n10241), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U11974 ( .A1(n10241), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U11975 ( .A1(n10241), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U11976 ( .A1(n10241), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U11977 ( .A1(n10241), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U11978 ( .A1(n10241), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U11979 ( .A1(n10241), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U11980 ( .A1(n10241), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U11981 ( .A1(n10241), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U11982 ( .A1(n10241), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U11983 ( .A1(n10241), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U11984 ( .A1(n10241), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U11985 ( .A1(n10241), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U11986 ( .A1(n10241), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U11987 ( .A1(n10241), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U11988 ( .A1(n10241), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  OAI21_X1 U11989 ( .B1(n10242), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10243) );
  XNOR2_X1 U11990 ( .A(n10243), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11863) );
  INV_X1 U11991 ( .A(n11863), .ZN(n10676) );
  INV_X1 U11992 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10244) );
  OAI222_X1 U11993 ( .A1(n10676), .A2(P1_U3086), .B1(n15990), .B2(n10245), 
        .C1(n10244), .C2(n15992), .ZN(P1_U3344) );
  INV_X1 U11994 ( .A(SI_13_), .ZN(n10247) );
  OAI222_X1 U11995 ( .A1(P3_U3151), .A2(n12498), .B1(n14150), .B2(n10247), 
        .C1(n14154), .C2(n10246), .ZN(P3_U3282) );
  INV_X1 U11996 ( .A(n11959), .ZN(n10253) );
  OAI222_X1 U11997 ( .A1(n15131), .A2(n10253), .B1(n16126), .B2(P2_U3088), 
        .C1(n10248), .C2(n15133), .ZN(P2_U3315) );
  NAND2_X1 U11998 ( .A1(n10250), .A2(n10249), .ZN(n10384) );
  NAND2_X1 U11999 ( .A1(n10384), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10251) );
  XNOR2_X1 U12000 ( .A(n10251), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11960) );
  INV_X1 U12001 ( .A(n11960), .ZN(n10836) );
  OAI222_X1 U12002 ( .A1(P1_U3086), .A2(n10836), .B1(n15990), .B2(n10253), 
        .C1(n10252), .C2(n15992), .ZN(P1_U3343) );
  XNOR2_X1 U12003 ( .A(n10372), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n10279) );
  MUX2_X1 U12004 ( .A(n8578), .B(P2_REG2_REG_1__SCAN_IN), .S(n16045), .Z(
        n16043) );
  AND2_X1 U12005 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n16042) );
  NAND2_X1 U12006 ( .A1(n16043), .A2(n16042), .ZN(n16041) );
  INV_X1 U12007 ( .A(n16045), .ZN(n10254) );
  NAND2_X1 U12008 ( .A1(n10254), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10255) );
  NAND2_X1 U12009 ( .A1(n16041), .A2(n10255), .ZN(n16054) );
  XNOR2_X1 U12010 ( .A(n10282), .B(n10256), .ZN(n16055) );
  NAND2_X1 U12011 ( .A1(n16054), .A2(n16055), .ZN(n16053) );
  NAND2_X1 U12012 ( .A1(n10282), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10257) );
  NAND2_X1 U12013 ( .A1(n16053), .A2(n10257), .ZN(n14739) );
  XNOR2_X1 U12014 ( .A(n14745), .B(n10258), .ZN(n14740) );
  NAND2_X1 U12015 ( .A1(n14739), .A2(n14740), .ZN(n14738) );
  NAND2_X1 U12016 ( .A1(n14745), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10259) );
  NAND2_X1 U12017 ( .A1(n14738), .A2(n10259), .ZN(n16066) );
  XNOR2_X1 U12018 ( .A(n10287), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n16067) );
  NAND2_X1 U12019 ( .A1(n16066), .A2(n16067), .ZN(n16065) );
  NAND2_X1 U12020 ( .A1(n16071), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10260) );
  NAND2_X1 U12021 ( .A1(n16065), .A2(n10260), .ZN(n14751) );
  INV_X1 U12022 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10261) );
  MUX2_X1 U12023 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10261), .S(n14756), .Z(
        n14752) );
  NAND2_X1 U12024 ( .A1(n14751), .A2(n14752), .ZN(n14750) );
  NAND2_X1 U12025 ( .A1(n14756), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10262) );
  NAND2_X1 U12026 ( .A1(n14750), .A2(n10262), .ZN(n14763) );
  XNOR2_X1 U12027 ( .A(n14769), .B(n11931), .ZN(n14764) );
  NAND2_X1 U12028 ( .A1(n14763), .A2(n14764), .ZN(n14762) );
  NAND2_X1 U12029 ( .A1(n14769), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10263) );
  NAND2_X1 U12030 ( .A1(n14762), .A2(n10263), .ZN(n14777) );
  XNOR2_X1 U12031 ( .A(n14783), .B(n10264), .ZN(n14778) );
  NAND2_X1 U12032 ( .A1(n14777), .A2(n14778), .ZN(n14776) );
  NAND2_X1 U12033 ( .A1(n14783), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10265) );
  NAND2_X1 U12034 ( .A1(n14776), .A2(n10265), .ZN(n14790) );
  INV_X1 U12035 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10266) );
  XNOR2_X1 U12036 ( .A(n14797), .B(n10266), .ZN(n14791) );
  NAND2_X1 U12037 ( .A1(n14790), .A2(n14791), .ZN(n16140) );
  XNOR2_X1 U12038 ( .A(n16151), .B(n12098), .ZN(n16142) );
  NAND2_X1 U12039 ( .A1(n14797), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n16139) );
  AND2_X1 U12040 ( .A1(n16142), .A2(n16139), .ZN(n10267) );
  NAND2_X1 U12041 ( .A1(n16140), .A2(n10267), .ZN(n16141) );
  NAND2_X1 U12042 ( .A1(n10304), .A2(n12098), .ZN(n10268) );
  NAND2_X1 U12043 ( .A1(n16141), .A2(n10268), .ZN(n10278) );
  OR2_X1 U12044 ( .A1(n10278), .A2(n10279), .ZN(n10364) );
  INV_X1 U12045 ( .A(n10364), .ZN(n10277) );
  NAND2_X1 U12046 ( .A1(n10270), .A2(n10269), .ZN(n10275) );
  OAI21_X1 U12047 ( .B1(n10273), .B2(n10272), .A(n10271), .ZN(n10274) );
  NAND2_X1 U12048 ( .A1(n10275), .A2(n10274), .ZN(n10312) );
  OR2_X1 U12049 ( .A1(n15115), .A2(P2_U3088), .ZN(n10276) );
  OR2_X1 U12050 ( .A1(n10312), .A2(n10276), .ZN(n10307) );
  AOI211_X1 U12051 ( .C1(n10279), .C2(n10278), .A(n10277), .B(n16114), .ZN(
        n10317) );
  MUX2_X1 U12052 ( .A(n10280), .B(P2_REG1_REG_1__SCAN_IN), .S(n16045), .Z(
        n16048) );
  AND2_X1 U12053 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n16049) );
  NAND2_X1 U12054 ( .A1(n16048), .A2(n16049), .ZN(n16047) );
  OAI21_X1 U12055 ( .B1(n10280), .B2(n16045), .A(n16047), .ZN(n16060) );
  INV_X1 U12056 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10281) );
  XNOR2_X1 U12057 ( .A(n10282), .B(n10281), .ZN(n16059) );
  NAND2_X1 U12058 ( .A1(n16060), .A2(n16059), .ZN(n10284) );
  NAND2_X1 U12059 ( .A1(n10282), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10283) );
  NAND2_X1 U12060 ( .A1(n10284), .A2(n10283), .ZN(n14742) );
  MUX2_X1 U12061 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10285), .S(n14745), .Z(
        n14743) );
  NAND2_X1 U12062 ( .A1(n14742), .A2(n14743), .ZN(n14741) );
  NAND2_X1 U12063 ( .A1(n14745), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10286) );
  NAND2_X1 U12064 ( .A1(n14741), .A2(n10286), .ZN(n16074) );
  INV_X1 U12065 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10288) );
  MUX2_X1 U12066 ( .A(n10288), .B(P2_REG1_REG_4__SCAN_IN), .S(n10287), .Z(
        n16073) );
  NAND2_X1 U12067 ( .A1(n16074), .A2(n16073), .ZN(n16072) );
  NAND2_X1 U12068 ( .A1(n16071), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n14754) );
  NAND2_X1 U12069 ( .A1(n16072), .A2(n14754), .ZN(n10291) );
  MUX2_X1 U12070 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10289), .S(n14756), .Z(
        n10290) );
  NAND2_X1 U12071 ( .A1(n10291), .A2(n10290), .ZN(n14767) );
  NAND2_X1 U12072 ( .A1(n14756), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n14766) );
  NAND2_X1 U12073 ( .A1(n14767), .A2(n14766), .ZN(n10294) );
  MUX2_X1 U12074 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10292), .S(n14769), .Z(
        n10293) );
  NAND2_X1 U12075 ( .A1(n10294), .A2(n10293), .ZN(n14781) );
  NAND2_X1 U12076 ( .A1(n14769), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n14780) );
  NAND2_X1 U12077 ( .A1(n14781), .A2(n14780), .ZN(n10297) );
  INV_X1 U12078 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10295) );
  MUX2_X1 U12079 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10295), .S(n14783), .Z(
        n10296) );
  NAND2_X1 U12080 ( .A1(n10297), .A2(n10296), .ZN(n14794) );
  NAND2_X1 U12081 ( .A1(n14783), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n14793) );
  NAND2_X1 U12082 ( .A1(n14794), .A2(n14793), .ZN(n10300) );
  MUX2_X1 U12083 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10298), .S(n14797), .Z(
        n10299) );
  NAND2_X1 U12084 ( .A1(n10300), .A2(n10299), .ZN(n14796) );
  NAND2_X1 U12085 ( .A1(n14797), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10301) );
  NAND2_X1 U12086 ( .A1(n14796), .A2(n10301), .ZN(n16144) );
  INV_X1 U12087 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10302) );
  MUX2_X1 U12088 ( .A(n10302), .B(P2_REG1_REG_9__SCAN_IN), .S(n16151), .Z(
        n10303) );
  OR2_X1 U12089 ( .A1(n16144), .A2(n10303), .ZN(n16145) );
  NAND2_X1 U12090 ( .A1(n10304), .A2(n10302), .ZN(n10305) );
  NAND2_X1 U12091 ( .A1(n16145), .A2(n10305), .ZN(n10310) );
  INV_X1 U12092 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n16576) );
  MUX2_X1 U12093 ( .A(n16576), .B(P2_REG1_REG_10__SCAN_IN), .S(n10372), .Z(
        n10309) );
  OR2_X1 U12094 ( .A1(n10310), .A2(n10309), .ZN(n10378) );
  INV_X1 U12095 ( .A(n10378), .ZN(n10308) );
  AOI211_X1 U12096 ( .C1(n10310), .C2(n10309), .A(n10308), .B(n11858), .ZN(
        n10316) );
  OR2_X1 U12097 ( .A1(n10312), .A2(n10311), .ZN(n16087) );
  AND2_X1 U12098 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11467) );
  AOI21_X1 U12099 ( .B1(n16110), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n11467), 
        .ZN(n10313) );
  OAI21_X1 U12100 ( .B1(n16127), .B2(n10314), .A(n10313), .ZN(n10315) );
  OR3_X1 U12101 ( .A1(n10317), .A2(n10316), .A3(n10315), .ZN(P2_U3224) );
  NAND2_X1 U12102 ( .A1(n10319), .A2(n10318), .ZN(n16164) );
  INV_X1 U12103 ( .A(n13373), .ZN(n10417) );
  OR2_X1 U12104 ( .A1(n16164), .A2(n10417), .ZN(n15511) );
  OR3_X1 U12105 ( .A1(n16164), .A2(n15982), .A3(n13373), .ZN(n15512) );
  XNOR2_X1 U12106 ( .A(n10471), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n15393) );
  AND2_X1 U12107 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n15392) );
  NAND2_X1 U12108 ( .A1(n15393), .A2(n15392), .ZN(n15391) );
  INV_X1 U12109 ( .A(n10471), .ZN(n15390) );
  NAND2_X1 U12110 ( .A1(n15390), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10320) );
  NAND2_X1 U12111 ( .A1(n15391), .A2(n10320), .ZN(n15402) );
  XNOR2_X1 U12112 ( .A(n15404), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n15401) );
  NAND2_X1 U12113 ( .A1(n15402), .A2(n15401), .ZN(n10323) );
  INV_X1 U12114 ( .A(n15404), .ZN(n10321) );
  NAND2_X1 U12115 ( .A1(n10321), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n10322) );
  NAND2_X1 U12116 ( .A1(n10323), .A2(n10322), .ZN(n15414) );
  INV_X1 U12117 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10505) );
  MUX2_X1 U12118 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10505), .S(n15412), .Z(
        n15415) );
  NAND2_X1 U12119 ( .A1(n15414), .A2(n15415), .ZN(n15413) );
  NAND2_X1 U12120 ( .A1(n15412), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n10327) );
  NAND2_X1 U12121 ( .A1(n15413), .A2(n10327), .ZN(n10325) );
  INV_X1 U12122 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10528) );
  MUX2_X1 U12123 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10528), .S(n10755), .Z(
        n10324) );
  NAND2_X1 U12124 ( .A1(n10325), .A2(n10324), .ZN(n15434) );
  MUX2_X1 U12125 ( .A(n10528), .B(P1_REG2_REG_4__SCAN_IN), .S(n10755), .Z(
        n10326) );
  NAND3_X1 U12126 ( .A1(n15413), .A2(n10327), .A3(n10326), .ZN(n10328) );
  AND3_X1 U12127 ( .A1(n15516), .A2(n15434), .A3(n10328), .ZN(n10335) );
  INV_X1 U12128 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n16208) );
  NAND2_X1 U12129 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n10775) );
  INV_X1 U12130 ( .A(n15982), .ZN(n16159) );
  INV_X1 U12131 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n16413) );
  MUX2_X1 U12132 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n16413), .S(n10471), .Z(
        n15387) );
  NAND2_X1 U12133 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n15388) );
  AOI21_X1 U12134 ( .B1(n15390), .B2(P1_REG1_REG_1__SCAN_IN), .A(n15386), .ZN(
        n15400) );
  INV_X1 U12135 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n16440) );
  MUX2_X1 U12136 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n16440), .S(n15404), .Z(
        n15399) );
  NOR2_X1 U12137 ( .A1(n15400), .A2(n15399), .ZN(n15418) );
  NOR2_X1 U12138 ( .A1(n15404), .A2(n16440), .ZN(n15417) );
  INV_X1 U12139 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10504) );
  MUX2_X1 U12140 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10504), .S(n15412), .Z(
        n15416) );
  OAI21_X1 U12141 ( .B1(n15418), .B2(n15417), .A(n15416), .ZN(n15420) );
  NAND2_X1 U12142 ( .A1(n15412), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10330) );
  INV_X1 U12143 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n16468) );
  MUX2_X1 U12144 ( .A(n16468), .B(P1_REG1_REG_4__SCAN_IN), .S(n10755), .Z(
        n10329) );
  INV_X1 U12145 ( .A(n10436), .ZN(n10332) );
  NAND3_X1 U12146 ( .A1(n15420), .A2(n10330), .A3(n10329), .ZN(n10331) );
  NAND3_X1 U12147 ( .A1(n15517), .A2(n10332), .A3(n10331), .ZN(n10333) );
  OAI211_X1 U12148 ( .C1(n15524), .C2(n16208), .A(n10775), .B(n10333), .ZN(
        n10334) );
  AOI211_X1 U12149 ( .C1(n15477), .C2(n10755), .A(n10335), .B(n10334), .ZN(
        n10362) );
  INV_X1 U12150 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n16401) );
  AOI21_X1 U12151 ( .B1(n16159), .B2(n16401), .A(n13373), .ZN(n16158) );
  NAND2_X1 U12152 ( .A1(n10336), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10337) );
  INV_X1 U12153 ( .A(n10410), .ZN(n10338) );
  INV_X1 U12154 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n16160) );
  NOR2_X1 U12155 ( .A1(n10468), .A2(n10339), .ZN(n10340) );
  XNOR2_X1 U12156 ( .A(n10340), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n15998) );
  MUX2_X1 U12157 ( .A(n16160), .B(n15998), .S(n13204), .Z(n13308) );
  INV_X1 U12158 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n16390) );
  OAI22_X1 U12159 ( .A1(n15136), .A2(n13308), .B1(n10410), .B2(n16390), .ZN(
        n10341) );
  INV_X1 U12160 ( .A(n10341), .ZN(n10356) );
  XNOR2_X2 U12161 ( .A(n10343), .B(n10342), .ZN(n15976) );
  INV_X1 U12162 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10344) );
  NAND2_X1 U12163 ( .A1(n13277), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10354) );
  INV_X1 U12164 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10349) );
  NAND2_X4 U12165 ( .A1(n10350), .A2(n15976), .ZN(n13284) );
  NAND2_X2 U12166 ( .A1(n15979), .A2(n15976), .ZN(n13279) );
  INV_X1 U12167 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10351) );
  OR2_X1 U12168 ( .A1(n13279), .A2(n10351), .ZN(n10352) );
  NAND2_X1 U12169 ( .A1(n15385), .A2(n7432), .ZN(n10355) );
  NAND2_X1 U12170 ( .A1(n10356), .A2(n10355), .ZN(n10465) );
  INV_X1 U12171 ( .A(n12984), .ZN(n12999) );
  NAND2_X1 U12172 ( .A1(n10357), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10358) );
  NAND2_X1 U12173 ( .A1(n16386), .A2(n10409), .ZN(n15810) );
  OAI22_X1 U12174 ( .A1(n7462), .A2(n13308), .B1(n10410), .B2(n16160), .ZN(
        n10359) );
  AOI21_X1 U12175 ( .B1(n15252), .B2(n15385), .A(n10359), .ZN(n10466) );
  XOR2_X1 U12176 ( .A(n10465), .B(n10466), .Z(n10429) );
  MUX2_X1 U12177 ( .A(n15392), .B(n10429), .S(n15982), .Z(n10360) );
  NAND2_X1 U12178 ( .A1(n10360), .A2(n10417), .ZN(n10361) );
  OAI211_X1 U12179 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n16158), .A(n10361), .B(
        P1_U4016), .ZN(n15409) );
  NAND2_X1 U12180 ( .A1(n10362), .A2(n15409), .ZN(P1_U3247) );
  XNOR2_X1 U12181 ( .A(n10576), .B(P2_REG2_REG_11__SCAN_IN), .ZN(n10367) );
  NAND2_X1 U12182 ( .A1(n10372), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10363) );
  NAND2_X1 U12183 ( .A1(n10364), .A2(n10363), .ZN(n10366) );
  OR2_X1 U12184 ( .A1(n10366), .A2(n10367), .ZN(n16132) );
  INV_X1 U12185 ( .A(n16132), .ZN(n10365) );
  AOI21_X1 U12186 ( .B1(n10367), .B2(n10366), .A(n10365), .ZN(n10382) );
  NOR2_X1 U12187 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10368), .ZN(n10371) );
  INV_X1 U12188 ( .A(n10576), .ZN(n10369) );
  NOR2_X1 U12189 ( .A1(n16127), .A2(n10369), .ZN(n10370) );
  AOI211_X1 U12190 ( .C1(n16110), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n10371), 
        .B(n10370), .ZN(n10381) );
  NAND2_X1 U12191 ( .A1(n10372), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10377) );
  NAND2_X1 U12192 ( .A1(n10378), .A2(n10377), .ZN(n10375) );
  INV_X1 U12193 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10373) );
  MUX2_X1 U12194 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10373), .S(n10576), .Z(
        n10374) );
  NAND2_X1 U12195 ( .A1(n10375), .A2(n10374), .ZN(n10568) );
  MUX2_X1 U12196 ( .A(n10373), .B(P2_REG1_REG_11__SCAN_IN), .S(n10576), .Z(
        n10376) );
  NAND3_X1 U12197 ( .A1(n10378), .A2(n10377), .A3(n10376), .ZN(n10379) );
  NAND3_X1 U12198 ( .A1(n16148), .A2(n10568), .A3(n10379), .ZN(n10380) );
  OAI211_X1 U12199 ( .C1(n10382), .C2(n16114), .A(n10381), .B(n10380), .ZN(
        P2_U3225) );
  INV_X1 U12200 ( .A(n13628), .ZN(n13618) );
  OAI222_X1 U12201 ( .A1(P3_U3151), .A2(n13618), .B1(n14150), .B2(n14435), 
        .C1(n14154), .C2(n10383), .ZN(P3_U3281) );
  NAND2_X1 U12202 ( .A1(n10387), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10386) );
  INV_X1 U12203 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10385) );
  MUX2_X1 U12204 ( .A(n10386), .B(P1_IR_REG_31__SCAN_IN), .S(n10385), .Z(
        n10388) );
  NAND2_X1 U12205 ( .A1(n10388), .A2(n10648), .ZN(n11445) );
  INV_X1 U12206 ( .A(n11999), .ZN(n10491) );
  OAI222_X1 U12207 ( .A1(P1_U3086), .A2(n11445), .B1(n15990), .B2(n10491), 
        .C1(n10389), .C2(n15992), .ZN(P1_U3342) );
  INV_X1 U12208 ( .A(n10401), .ZN(n10392) );
  NOR2_X1 U12209 ( .A1(n10424), .A2(n11053), .ZN(n10406) );
  NAND2_X1 U12210 ( .A1(n15985), .A2(n15991), .ZN(n15968) );
  OAI21_X1 U12211 ( .B1(n10392), .B2(P1_D_REG_1__SCAN_IN), .A(n15968), .ZN(
        n10858) );
  INV_X1 U12212 ( .A(n10858), .ZN(n10404) );
  NOR4_X1 U12213 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n10396) );
  NOR4_X1 U12214 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n10395) );
  NOR4_X1 U12215 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n10394) );
  NOR4_X1 U12216 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n10393) );
  NAND4_X1 U12217 ( .A1(n10396), .A2(n10395), .A3(n10394), .A4(n10393), .ZN(
        n10403) );
  NOR2_X1 U12218 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n10400) );
  NOR4_X1 U12219 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n10399) );
  NOR4_X1 U12220 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n10398) );
  NOR4_X1 U12221 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n10397) );
  NAND4_X1 U12222 ( .A1(n10400), .A2(n10399), .A3(n10398), .A4(n10397), .ZN(
        n10402) );
  OAI21_X1 U12223 ( .B1(n10403), .B2(n10402), .A(n10401), .ZN(n10857) );
  NAND2_X1 U12224 ( .A1(n10404), .A2(n10857), .ZN(n11119) );
  INV_X1 U12225 ( .A(n11119), .ZN(n10405) );
  NAND2_X1 U12226 ( .A1(n10406), .A2(n10405), .ZN(n10423) );
  INV_X1 U12227 ( .A(n16386), .ZN(n10407) );
  NAND2_X1 U12228 ( .A1(n16556), .A2(n12995), .ZN(n10408) );
  OR2_X1 U12229 ( .A1(n12995), .A2(n10409), .ZN(n10415) );
  NAND3_X1 U12230 ( .A1(n10415), .A2(n10411), .A3(n10410), .ZN(n10856) );
  INV_X1 U12231 ( .A(n10856), .ZN(n10414) );
  NAND2_X1 U12232 ( .A1(n12993), .A2(n13341), .ZN(n16392) );
  INV_X1 U12233 ( .A(n16392), .ZN(n10412) );
  NAND2_X1 U12234 ( .A1(n12983), .A2(n10412), .ZN(n16493) );
  OAI21_X1 U12235 ( .B1(n11119), .B2(n11053), .A(n10859), .ZN(n10413) );
  NAND2_X1 U12236 ( .A1(n10414), .A2(n10413), .ZN(n10527) );
  NOR2_X1 U12237 ( .A1(n10527), .A2(P1_U3086), .ZN(n10515) );
  INV_X1 U12238 ( .A(n10515), .ZN(n10427) );
  INV_X1 U12239 ( .A(n10415), .ZN(n10416) );
  INV_X1 U12240 ( .A(n15264), .ZN(n15277) );
  NAND2_X1 U12241 ( .A1(n15277), .A2(n15789), .ZN(n15362) );
  INV_X4 U12242 ( .A(n13279), .ZN(n13170) );
  NAND2_X1 U12243 ( .A1(n13170), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n10421) );
  INV_X1 U12244 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n11129) );
  OR2_X1 U12245 ( .A1(n10529), .A2(n11129), .ZN(n10420) );
  INV_X1 U12246 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n11130) );
  OR2_X1 U12247 ( .A1(n10797), .A2(n11130), .ZN(n10418) );
  NAND4_X4 U12248 ( .A1(n10421), .A2(n10420), .A3(n10419), .A4(n10418), .ZN(
        n15384) );
  INV_X1 U12249 ( .A(n12993), .ZN(n12998) );
  AND2_X1 U12250 ( .A1(n16386), .A2(n12998), .ZN(n11128) );
  INV_X1 U12251 ( .A(n11128), .ZN(n10422) );
  OR2_X1 U12252 ( .A1(n10423), .A2(n10422), .ZN(n10425) );
  OAI22_X1 U12253 ( .A1(n15362), .A2(n7600), .B1(n15340), .B2(n13308), .ZN(
        n10426) );
  AOI21_X1 U12254 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n10427), .A(n10426), .ZN(
        n10428) );
  OAI21_X1 U12255 ( .B1(n15367), .B2(n10429), .A(n10428), .ZN(P1_U3232) );
  NAND2_X1 U12256 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n10908) );
  NAND2_X1 U12257 ( .A1(n10755), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n15433) );
  NAND2_X1 U12258 ( .A1(n15434), .A2(n15433), .ZN(n10431) );
  INV_X1 U12259 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10769) );
  MUX2_X1 U12260 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10769), .S(n15431), .Z(
        n10430) );
  NAND2_X1 U12261 ( .A1(n10431), .A2(n10430), .ZN(n15436) );
  NAND2_X1 U12262 ( .A1(n15431), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10432) );
  NAND2_X1 U12263 ( .A1(n15436), .A2(n10432), .ZN(n10434) );
  INV_X1 U12264 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11210) );
  MUX2_X1 U12265 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11210), .S(n10893), .Z(
        n10433) );
  NAND2_X1 U12266 ( .A1(n10434), .A2(n10433), .ZN(n15446) );
  OAI211_X1 U12267 ( .C1(n10434), .C2(n10433), .A(n15516), .B(n15446), .ZN(
        n10435) );
  NAND2_X1 U12268 ( .A1(n10908), .A2(n10435), .ZN(n10442) );
  AOI21_X1 U12269 ( .B1(n10755), .B2(P1_REG1_REG_4__SCAN_IN), .A(n10436), .ZN(
        n15428) );
  INV_X1 U12270 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10437) );
  MUX2_X1 U12271 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10437), .S(n15431), .Z(
        n15429) );
  NAND2_X1 U12272 ( .A1(n15428), .A2(n15429), .ZN(n15427) );
  OAI21_X1 U12273 ( .B1(n15431), .B2(P1_REG1_REG_5__SCAN_IN), .A(n15427), .ZN(
        n10440) );
  INV_X1 U12274 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n16496) );
  MUX2_X1 U12275 ( .A(n16496), .B(P1_REG1_REG_6__SCAN_IN), .S(n10893), .Z(
        n10439) );
  OR2_X1 U12276 ( .A1(n10440), .A2(n10439), .ZN(n15451) );
  INV_X1 U12277 ( .A(n15451), .ZN(n10438) );
  AOI211_X1 U12278 ( .C1(n10440), .C2(n10439), .A(n15398), .B(n10438), .ZN(
        n10441) );
  AOI211_X1 U12279 ( .C1(n16162), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n10442), .B(
        n10441), .ZN(n10443) );
  OAI21_X1 U12280 ( .B1(n10444), .B2(n15511), .A(n10443), .ZN(P1_U3249) );
  NOR2_X1 U12281 ( .A1(n10446), .A2(n10445), .ZN(n11318) );
  AND2_X1 U12282 ( .A1(n16040), .A2(n11315), .ZN(n16032) );
  INV_X1 U12283 ( .A(n16039), .ZN(n10448) );
  XNOR2_X1 U12284 ( .A(n10605), .B(n10604), .ZN(n11793) );
  XNOR2_X1 U12285 ( .A(n11319), .B(n9157), .ZN(n10449) );
  INV_X1 U12286 ( .A(n10450), .ZN(n16610) );
  INV_X1 U12287 ( .A(n10716), .ZN(n11791) );
  INV_X1 U12288 ( .A(n16420), .ZN(n10451) );
  NAND2_X1 U12289 ( .A1(n10451), .A2(n10660), .ZN(n10620) );
  NAND2_X1 U12290 ( .A1(n10716), .A2(n10620), .ZN(n10452) );
  NAND2_X1 U12291 ( .A1(n10452), .A2(n14930), .ZN(n10453) );
  OR2_X1 U12292 ( .A1(n10453), .A2(n10608), .ZN(n11788) );
  OAI21_X1 U12293 ( .B1(n11791), .B2(n16616), .A(n11788), .ZN(n10454) );
  AOI21_X1 U12294 ( .B1(n11793), .B2(n16621), .A(n10454), .ZN(n10463) );
  INV_X1 U12295 ( .A(n10659), .ZN(n10623) );
  NAND2_X1 U12296 ( .A1(n10622), .A2(n10623), .ZN(n10456) );
  INV_X1 U12297 ( .A(n14735), .ZN(n10665) );
  NAND2_X1 U12298 ( .A1(n10665), .A2(n16420), .ZN(n10455) );
  NAND2_X1 U12299 ( .A1(n10456), .A2(n10455), .ZN(n10611) );
  XNOR2_X1 U12300 ( .A(n10611), .B(n10610), .ZN(n10462) );
  OR2_X1 U12301 ( .A1(n9155), .A2(n12139), .ZN(n10458) );
  NAND2_X1 U12302 ( .A1(n8519), .A2(n11851), .ZN(n10457) );
  NAND2_X1 U12303 ( .A1(n14733), .A2(n14913), .ZN(n10460) );
  NAND2_X1 U12304 ( .A1(n14735), .A2(n14911), .ZN(n10459) );
  AND2_X1 U12305 ( .A1(n10460), .A2(n10459), .ZN(n10707) );
  INV_X1 U12306 ( .A(n10707), .ZN(n10461) );
  AOI21_X1 U12307 ( .B1(n10462), .B2(n14981), .A(n10461), .ZN(n11795) );
  AND2_X1 U12308 ( .A1(n10463), .A2(n11795), .ZN(n16443) );
  NAND2_X1 U12309 ( .A1(n16622), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10464) );
  OAI21_X1 U12310 ( .B1(n16622), .B2(n16443), .A(n10464), .ZN(P2_U3501) );
  INV_X2 U12311 ( .A(n15221), .ZN(n15253) );
  MUX2_X1 U12312 ( .A(n15253), .B(n10466), .S(n10465), .Z(n10482) );
  NAND2_X1 U12313 ( .A1(n15384), .A2(n7432), .ZN(n10473) );
  OR2_X1 U12314 ( .A1(n12973), .A2(n10467), .ZN(n10470) );
  OR2_X1 U12315 ( .A1(n15136), .A2(n7601), .ZN(n10472) );
  NAND2_X1 U12316 ( .A1(n10473), .A2(n10472), .ZN(n10474) );
  NOR2_X1 U12317 ( .A1(n7601), .A2(n7462), .ZN(n10475) );
  AOI21_X1 U12318 ( .B1(n15252), .B2(n15384), .A(n10475), .ZN(n10477) );
  NAND2_X1 U12319 ( .A1(n10476), .A2(n10477), .ZN(n10499) );
  INV_X1 U12320 ( .A(n10476), .ZN(n10479) );
  INV_X1 U12321 ( .A(n10477), .ZN(n10478) );
  NAND2_X1 U12322 ( .A1(n10479), .A2(n10478), .ZN(n10480) );
  AND2_X1 U12323 ( .A1(n10499), .A2(n10480), .ZN(n10481) );
  NAND2_X1 U12324 ( .A1(n10481), .A2(n10482), .ZN(n10500) );
  OAI21_X1 U12325 ( .B1(n10482), .B2(n10481), .A(n10500), .ZN(n10489) );
  NAND2_X1 U12326 ( .A1(n13170), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n10486) );
  INV_X1 U12327 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10514) );
  OR2_X1 U12328 ( .A1(n10529), .A2(n10514), .ZN(n10485) );
  INV_X1 U12329 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n11141) );
  OR2_X1 U12330 ( .A1(n10797), .A2(n11141), .ZN(n10483) );
  OAI22_X1 U12331 ( .A1(n15362), .A2(n7856), .B1(n10515), .B2(n11129), .ZN(
        n10488) );
  NAND2_X1 U12332 ( .A1(n15277), .A2(n15787), .ZN(n15359) );
  INV_X1 U12333 ( .A(n15385), .ZN(n11123) );
  OAI22_X1 U12334 ( .A1(n15359), .A2(n11123), .B1(n15340), .B2(n7601), .ZN(
        n10487) );
  AOI211_X1 U12335 ( .C1(n15332), .C2(n10489), .A(n10488), .B(n10487), .ZN(
        n10490) );
  INV_X1 U12336 ( .A(n10490), .ZN(P1_U3222) );
  INV_X1 U12337 ( .A(n10572), .ZN(n10690) );
  OAI222_X1 U12338 ( .A1(n15133), .A2(n10492), .B1(n10690), .B2(P2_U3088), 
        .C1(n15123), .C2(n10491), .ZN(P2_U3314) );
  NAND2_X1 U12339 ( .A1(n15383), .A2(n7432), .ZN(n10495) );
  OAI21_X1 U12340 ( .B1(n16434), .B2(n15136), .A(n10495), .ZN(n10496) );
  XNOR2_X1 U12341 ( .A(n10496), .B(n15221), .ZN(n10524) );
  OR2_X1 U12342 ( .A1(n16434), .A2(n7462), .ZN(n10497) );
  NAND2_X1 U12343 ( .A1(n10498), .A2(n10497), .ZN(n10522) );
  XNOR2_X1 U12344 ( .A(n10524), .B(n10522), .ZN(n10502) );
  NAND2_X1 U12345 ( .A1(n10500), .A2(n10499), .ZN(n10501) );
  NAND2_X1 U12346 ( .A1(n10501), .A2(n10502), .ZN(n10525) );
  OAI21_X1 U12347 ( .B1(n10502), .B2(n10501), .A(n10525), .ZN(n10503) );
  NAND2_X1 U12348 ( .A1(n10503), .A2(n15332), .ZN(n10513) );
  NAND2_X1 U12349 ( .A1(n13170), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n10509) );
  OR2_X1 U12350 ( .A1(n10529), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10508) );
  OR2_X1 U12351 ( .A1(n13284), .A2(n10504), .ZN(n10507) );
  OR2_X1 U12352 ( .A1(n10797), .A2(n10505), .ZN(n10506) );
  OR2_X1 U12353 ( .A1(n10876), .A2(n16389), .ZN(n10511) );
  NAND2_X1 U12354 ( .A1(n15787), .A2(n15384), .ZN(n10510) );
  NAND2_X1 U12355 ( .A1(n10511), .A2(n10510), .ZN(n16431) );
  AOI22_X1 U12356 ( .A1(n15277), .A2(n16431), .B1(n15365), .B2(n7857), .ZN(
        n10512) );
  OAI211_X1 U12357 ( .C1(n10515), .C2(n10514), .A(n10513), .B(n10512), .ZN(
        P1_U3237) );
  NAND2_X1 U12358 ( .A1(n10516), .A2(n13289), .ZN(n10517) );
  NAND2_X1 U12359 ( .A1(n11173), .A2(n15255), .ZN(n10518) );
  OAI21_X1 U12360 ( .B1(n10876), .B2(n7462), .A(n10518), .ZN(n10519) );
  XNOR2_X1 U12361 ( .A(n10519), .B(n15221), .ZN(n10751) );
  NAND2_X1 U12362 ( .A1(n11173), .A2(n7432), .ZN(n10520) );
  NAND2_X1 U12363 ( .A1(n10521), .A2(n10520), .ZN(n10752) );
  INV_X1 U12364 ( .A(n10522), .ZN(n10523) );
  NAND2_X1 U12365 ( .A1(n10524), .A2(n10523), .ZN(n10526) );
  NAND2_X1 U12366 ( .A1(n10765), .A2(n15332), .ZN(n10543) );
  INV_X1 U12367 ( .A(n15360), .ZN(n15312) );
  INV_X1 U12368 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n15410) );
  NAND2_X1 U12369 ( .A1(n13170), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n10536) );
  OR2_X1 U12370 ( .A1(n13256), .A2(n10528), .ZN(n10535) );
  INV_X1 U12371 ( .A(n10770), .ZN(n10532) );
  INV_X1 U12372 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10530) );
  NAND2_X1 U12373 ( .A1(n15410), .A2(n10530), .ZN(n10531) );
  NAND2_X1 U12374 ( .A1(n10532), .A2(n10531), .ZN(n11367) );
  OR2_X1 U12375 ( .A1(n13282), .A2(n11367), .ZN(n10534) );
  OR2_X1 U12376 ( .A1(n13284), .A2(n16468), .ZN(n10533) );
  OR2_X1 U12377 ( .A1(n10878), .A2(n16389), .ZN(n10538) );
  NAND2_X1 U12378 ( .A1(n15787), .A2(n15383), .ZN(n10537) );
  AND2_X1 U12379 ( .A1(n10538), .A2(n10537), .ZN(n16450) );
  INV_X1 U12380 ( .A(n16450), .ZN(n11176) );
  AOI22_X1 U12381 ( .A1(n15277), .A2(n11176), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10539) );
  OAI21_X1 U12382 ( .B1(n16452), .B2(n15340), .A(n10539), .ZN(n10540) );
  AOI21_X1 U12383 ( .B1(n15312), .B2(n15410), .A(n10540), .ZN(n10541) );
  OAI21_X1 U12384 ( .B1(n10543), .B2(n10542), .A(n10541), .ZN(P1_U3218) );
  INV_X1 U12385 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11600) );
  MUX2_X1 U12386 ( .A(n11600), .B(P1_REG1_REG_11__SCAN_IN), .S(n11863), .Z(
        n10547) );
  INV_X1 U12387 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n16566) );
  INV_X1 U12388 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n11823) );
  NAND2_X1 U12389 ( .A1(n10893), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n15450) );
  INV_X1 U12390 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n11082) );
  MUX2_X1 U12391 ( .A(n11082), .B(P1_REG1_REG_7__SCAN_IN), .S(n15443), .Z(
        n15449) );
  AOI21_X1 U12392 ( .B1(n15443), .B2(P1_REG1_REG_7__SCAN_IN), .A(n15448), .ZN(
        n15457) );
  INV_X1 U12393 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n11581) );
  MUX2_X1 U12394 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n11581), .S(n15462), .Z(
        n15458) );
  NAND2_X1 U12395 ( .A1(n15457), .A2(n15458), .ZN(n15472) );
  NAND2_X1 U12396 ( .A1(n10544), .A2(n11581), .ZN(n15470) );
  MUX2_X1 U12397 ( .A(n11823), .B(P1_REG1_REG_9__SCAN_IN), .S(n15478), .Z(
        n15471) );
  AOI21_X1 U12398 ( .B1(n15472), .B2(n15470), .A(n15471), .ZN(n15474) );
  MUX2_X1 U12399 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n16566), .S(n15492), .Z(
        n15487) );
  NAND2_X1 U12400 ( .A1(n15488), .A2(n15487), .ZN(n15486) );
  OAI21_X1 U12401 ( .B1(n16566), .B2(n15489), .A(n15486), .ZN(n10546) );
  NOR2_X1 U12402 ( .A1(n10546), .A2(n10547), .ZN(n10675) );
  AOI21_X1 U12403 ( .B1(n10547), .B2(n10546), .A(n10675), .ZN(n10565) );
  NAND2_X1 U12404 ( .A1(n10893), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n15445) );
  NAND2_X1 U12405 ( .A1(n15446), .A2(n15445), .ZN(n10549) );
  INV_X1 U12406 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11331) );
  MUX2_X1 U12407 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n11331), .S(n15443), .Z(
        n10548) );
  NAND2_X1 U12408 ( .A1(n10549), .A2(n10548), .ZN(n15465) );
  NAND2_X1 U12409 ( .A1(n15443), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n15464) );
  NAND2_X1 U12410 ( .A1(n15465), .A2(n15464), .ZN(n10551) );
  INV_X1 U12411 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11069) );
  MUX2_X1 U12412 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11069), .S(n15462), .Z(
        n10550) );
  NAND2_X1 U12413 ( .A1(n10551), .A2(n10550), .ZN(n15481) );
  NAND2_X1 U12414 ( .A1(n15462), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n15480) );
  NAND2_X1 U12415 ( .A1(n15481), .A2(n15480), .ZN(n10553) );
  INV_X1 U12416 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11303) );
  MUX2_X1 U12417 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11303), .S(n15478), .Z(
        n10552) );
  NAND2_X1 U12418 ( .A1(n10553), .A2(n10552), .ZN(n15495) );
  NAND2_X1 U12419 ( .A1(n15478), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n15494) );
  NAND2_X1 U12420 ( .A1(n15495), .A2(n15494), .ZN(n10555) );
  INV_X1 U12421 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11595) );
  MUX2_X1 U12422 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11595), .S(n15492), .Z(
        n10554) );
  NAND2_X1 U12423 ( .A1(n10555), .A2(n10554), .ZN(n15497) );
  NAND2_X1 U12424 ( .A1(n15492), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10558) );
  INV_X1 U12425 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10556) );
  MUX2_X1 U12426 ( .A(n10556), .B(P1_REG2_REG_11__SCAN_IN), .S(n11863), .Z(
        n10557) );
  AOI21_X1 U12427 ( .B1(n15497), .B2(n10558), .A(n10557), .ZN(n10678) );
  NAND3_X1 U12428 ( .A1(n15497), .A2(n10558), .A3(n10557), .ZN(n10559) );
  NAND2_X1 U12429 ( .A1(n15516), .A2(n10559), .ZN(n10560) );
  OR2_X1 U12430 ( .A1(n10678), .A2(n10560), .ZN(n10562) );
  AND2_X1 U12431 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n12059) );
  AOI21_X1 U12432 ( .B1(n16162), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n12059), 
        .ZN(n10561) );
  OAI211_X1 U12433 ( .C1(n15511), .C2(n10676), .A(n10562), .B(n10561), .ZN(
        n10563) );
  INV_X1 U12434 ( .A(n10563), .ZN(n10564) );
  OAI21_X1 U12435 ( .B1(n10565), .B2(n15398), .A(n10564), .ZN(P1_U3254) );
  INV_X1 U12436 ( .A(n12312), .ZN(n10602) );
  AOI22_X1 U12437 ( .A1(n11837), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n11163), .ZN(n10566) );
  OAI21_X1 U12438 ( .B1(n10602), .B2(n15131), .A(n10566), .ZN(P2_U3313) );
  NAND2_X1 U12439 ( .A1(n10576), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10567) );
  NAND2_X1 U12440 ( .A1(n10568), .A2(n10567), .ZN(n16123) );
  MUX2_X1 U12441 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n10569), .S(n16126), .Z(
        n16122) );
  NAND2_X1 U12442 ( .A1(n16126), .A2(n10569), .ZN(n10570) );
  NAND2_X1 U12443 ( .A1(n16125), .A2(n10570), .ZN(n10574) );
  NAND2_X1 U12444 ( .A1(n10572), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10693) );
  OAI21_X1 U12445 ( .B1(n10572), .B2(P2_REG1_REG_13__SCAN_IN), .A(n10693), 
        .ZN(n10571) );
  NOR2_X1 U12446 ( .A1(n10574), .A2(n10571), .ZN(n10700) );
  INV_X1 U12447 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n12432) );
  OR2_X1 U12448 ( .A1(n10572), .A2(n12432), .ZN(n10573) );
  OAI211_X1 U12449 ( .C1(P2_REG1_REG_13__SCAN_IN), .C2(n10690), .A(n10574), 
        .B(n10573), .ZN(n10575) );
  NAND2_X1 U12450 ( .A1(n10575), .A2(n16148), .ZN(n10583) );
  INV_X1 U12451 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n12203) );
  OR2_X1 U12452 ( .A1(n10576), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n16131) );
  MUX2_X1 U12453 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n12203), .S(n16126), .Z(
        n16130) );
  AOI21_X1 U12454 ( .B1(n16132), .B2(n16131), .A(n16130), .ZN(n16134) );
  AOI21_X1 U12455 ( .B1(n12203), .B2(n16126), .A(n16134), .ZN(n10578) );
  XNOR2_X1 U12456 ( .A(n10690), .B(P2_REG2_REG_13__SCAN_IN), .ZN(n10577) );
  NAND2_X1 U12457 ( .A1(n10578), .A2(n10577), .ZN(n10689) );
  OAI211_X1 U12458 ( .C1(n10578), .C2(n10577), .A(n10689), .B(n16152), .ZN(
        n10582) );
  NAND2_X1 U12459 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n12090)
         );
  INV_X1 U12460 ( .A(n12090), .ZN(n10580) );
  NOR2_X1 U12461 ( .A1(n16127), .A2(n10690), .ZN(n10579) );
  AOI211_X1 U12462 ( .C1(n16110), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n10580), 
        .B(n10579), .ZN(n10581) );
  OAI211_X1 U12463 ( .C1(n10700), .C2(n10583), .A(n10582), .B(n10581), .ZN(
        P2_U3227) );
  NOR2_X1 U12464 ( .A1(n16507), .A2(n14981), .ZN(n10584) );
  OAI22_X1 U12465 ( .A1(n11328), .A2(n10584), .B1(n10665), .B2(n14953), .ZN(
        n11322) );
  INV_X1 U12466 ( .A(n11322), .ZN(n10586) );
  INV_X1 U12467 ( .A(n11324), .ZN(n10585) );
  OAI211_X1 U12468 ( .C1(n11328), .C2(n10450), .A(n10586), .B(n10585), .ZN(
        n10631) );
  NAND2_X1 U12469 ( .A1(n7433), .A2(n10631), .ZN(n10587) );
  OAI21_X1 U12470 ( .B1(n7433), .B2(n10590), .A(n10587), .ZN(P2_U3499) );
  NAND2_X1 U12471 ( .A1(n16148), .A2(n10590), .ZN(n10588) );
  OAI211_X1 U12472 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n16114), .A(n10588), .B(
        n16127), .ZN(n10593) );
  OAI22_X1 U12473 ( .A1(n10590), .A2(n11858), .B1(n16114), .B2(n10589), .ZN(
        n10592) );
  MUX2_X1 U12474 ( .A(n10593), .B(n10592), .S(n10591), .Z(n10597) );
  INV_X1 U12475 ( .A(n16110), .ZN(n16156) );
  INV_X1 U12476 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10595) );
  OAI22_X1 U12477 ( .A1(n16156), .A2(n10595), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10594), .ZN(n10596) );
  OR2_X1 U12478 ( .A1(n10597), .A2(n10596), .ZN(P2_U3214) );
  INV_X1 U12479 ( .A(n10598), .ZN(n10599) );
  OAI222_X1 U12480 ( .A1(n14150), .A2(n14430), .B1(n14154), .B2(n10599), .C1(
        n16366), .C2(P3_U3151), .ZN(P3_U3280) );
  NAND2_X1 U12481 ( .A1(n10648), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10600) );
  XNOR2_X1 U12482 ( .A(n10600), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12313) );
  INV_X1 U12483 ( .A(n12313), .ZN(n11458) );
  OAI222_X1 U12484 ( .A1(n11458), .A2(P1_U3086), .B1(n15990), .B2(n10602), 
        .C1(n10601), .C2(n15992), .ZN(P1_U3341) );
  INV_X2 U12485 ( .A(n16623), .ZN(n15102) );
  INV_X1 U12486 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10617) );
  NAND2_X1 U12487 ( .A1(n10605), .A2(n10604), .ZN(n10607) );
  INV_X1 U12488 ( .A(n14734), .ZN(n10624) );
  NAND2_X1 U12489 ( .A1(n11791), .A2(n10624), .ZN(n10606) );
  NAND2_X1 U12490 ( .A1(n10607), .A2(n10606), .ZN(n10812) );
  INV_X1 U12491 ( .A(n10815), .ZN(n10811) );
  XNOR2_X1 U12492 ( .A(n10812), .B(n10811), .ZN(n11993) );
  NAND2_X1 U12493 ( .A1(n10608), .A2(n11990), .ZN(n10823) );
  OAI211_X1 U12494 ( .C1(n10608), .C2(n11990), .A(n14930), .B(n10823), .ZN(
        n11989) );
  OAI21_X1 U12495 ( .B1(n11990), .B2(n16616), .A(n11989), .ZN(n10609) );
  AOI21_X1 U12496 ( .B1(n11993), .B2(n16621), .A(n10609), .ZN(n10615) );
  NAND2_X1 U12497 ( .A1(n10611), .A2(n10610), .ZN(n10613) );
  NAND2_X1 U12498 ( .A1(n10624), .A2(n10716), .ZN(n10612) );
  NAND2_X1 U12499 ( .A1(n10613), .A2(n10612), .ZN(n10816) );
  XNOR2_X1 U12500 ( .A(n10815), .B(n10816), .ZN(n10614) );
  INV_X1 U12501 ( .A(n14732), .ZN(n10997) );
  OAI22_X1 U12502 ( .A1(n10624), .A2(n14951), .B1(n10997), .B2(n14953), .ZN(
        n14171) );
  AOI21_X1 U12503 ( .B1(n10614), .B2(n14981), .A(n14171), .ZN(n11996) );
  NAND2_X1 U12504 ( .A1(n10615), .A2(n11996), .ZN(n10618) );
  NAND2_X1 U12505 ( .A1(n10618), .A2(n15102), .ZN(n10616) );
  OAI21_X1 U12506 ( .B1(n15102), .B2(n10617), .A(n10616), .ZN(P2_U3439) );
  NAND2_X1 U12507 ( .A1(n10618), .A2(n7433), .ZN(n10619) );
  OAI21_X1 U12508 ( .B1(n7433), .B2(n10285), .A(n10619), .ZN(P2_U3502) );
  INV_X1 U12509 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10630) );
  XNOR2_X1 U12510 ( .A(n10622), .B(n14202), .ZN(n16416) );
  INV_X1 U12511 ( .A(n16416), .ZN(n10628) );
  INV_X1 U12512 ( .A(n10620), .ZN(n10621) );
  AOI211_X1 U12513 ( .C1(n8032), .C2(n16420), .A(n14986), .B(n10621), .ZN(
        n16418) );
  AOI21_X1 U12514 ( .B1(n15079), .B2(n16420), .A(n16418), .ZN(n10627) );
  XNOR2_X1 U12515 ( .A(n10623), .B(n10622), .ZN(n10626) );
  OAI22_X1 U12516 ( .A1(n10625), .A2(n14951), .B1(n10624), .B2(n14953), .ZN(
        n14204) );
  AOI21_X1 U12517 ( .B1(n10626), .B2(n14981), .A(n14204), .ZN(n16423) );
  OAI211_X1 U12518 ( .C1(n15082), .C2(n10628), .A(n10627), .B(n16423), .ZN(
        n15085) );
  NAND2_X1 U12519 ( .A1(n15102), .A2(n15085), .ZN(n10629) );
  OAI21_X1 U12520 ( .B1(n15102), .B2(n10630), .A(n10629), .ZN(P2_U3433) );
  INV_X1 U12521 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10633) );
  NAND2_X1 U12522 ( .A1(n15102), .A2(n10631), .ZN(n10632) );
  OAI21_X1 U12523 ( .B1(n15102), .B2(n10633), .A(n10632), .ZN(P2_U3430) );
  INV_X1 U12524 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n10635) );
  NAND2_X1 U12525 ( .A1(n12163), .A2(n11644), .ZN(n10634) );
  OAI21_X1 U12526 ( .B1(n11644), .B2(n10635), .A(n10634), .ZN(P3_U3496) );
  INV_X1 U12527 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n10638) );
  NAND2_X1 U12528 ( .A1(n10636), .A2(n11644), .ZN(n10637) );
  OAI21_X1 U12529 ( .B1(n11644), .B2(n10638), .A(n10637), .ZN(P3_U3491) );
  INV_X1 U12530 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n10640) );
  NAND2_X1 U12531 ( .A1(n13485), .A2(n11644), .ZN(n10639) );
  OAI21_X1 U12532 ( .B1(n11644), .B2(n10640), .A(n10639), .ZN(P3_U3495) );
  INV_X1 U12533 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n10642) );
  NAND2_X1 U12534 ( .A1(n12832), .A2(n11644), .ZN(n10641) );
  OAI21_X1 U12535 ( .B1(n11644), .B2(n10642), .A(n10641), .ZN(P3_U3501) );
  INV_X1 U12536 ( .A(n12402), .ZN(n10651) );
  INV_X1 U12537 ( .A(n16079), .ZN(n11842) );
  OAI222_X1 U12538 ( .A1(n15131), .A2(n10651), .B1(n11842), .B2(P2_U3088), 
        .C1(n10643), .C2(n15133), .ZN(P2_U3312) );
  INV_X1 U12539 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n10647) );
  INV_X1 U12540 ( .A(n10645), .ZN(n13483) );
  NAND2_X1 U12541 ( .A1(n13483), .A2(n11644), .ZN(n10646) );
  OAI21_X1 U12542 ( .B1(n11644), .B2(n10647), .A(n10646), .ZN(P3_U3493) );
  OAI21_X1 U12543 ( .B1(n10648), .B2(P1_IR_REG_14__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10649) );
  XNOR2_X1 U12544 ( .A(n10649), .B(P1_IR_REG_15__SCAN_IN), .ZN(n12403) );
  INV_X1 U12545 ( .A(n12403), .ZN(n12213) );
  OAI222_X1 U12546 ( .A1(P1_U3086), .A2(n12213), .B1(n15990), .B2(n10651), 
        .C1(n10650), .C2(n15992), .ZN(P1_U3340) );
  INV_X1 U12547 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n10653) );
  NAND2_X1 U12548 ( .A1(n13834), .A2(n11644), .ZN(n10652) );
  OAI21_X1 U12549 ( .B1(P3_U3897), .B2(n10653), .A(n10652), .ZN(P3_U3511) );
  INV_X1 U12550 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n10655) );
  NAND2_X1 U12551 ( .A1(n12394), .A2(n11644), .ZN(n10654) );
  OAI21_X1 U12552 ( .B1(n11644), .B2(n10655), .A(n10654), .ZN(P3_U3498) );
  INV_X1 U12553 ( .A(n10656), .ZN(n10657) );
  OAI222_X1 U12554 ( .A1(P3_U3151), .A2(n13649), .B1(n14150), .B2(n14429), 
        .C1(n14154), .C2(n10657), .ZN(P3_U3279) );
  INV_X1 U12555 ( .A(n14702), .ZN(n11464) );
  NAND2_X1 U12556 ( .A1(n14707), .A2(n14884), .ZN(n14694) );
  INV_X1 U12557 ( .A(n14694), .ZN(n14671) );
  NAND2_X1 U12558 ( .A1(n14671), .A2(n14737), .ZN(n10658) );
  MUX2_X1 U12559 ( .A(n10658), .B(n14705), .S(n8032), .Z(n10664) );
  OAI21_X1 U12560 ( .B1(n10660), .B2(n14884), .A(n10659), .ZN(n10662) );
  OR2_X1 U12561 ( .A1(n10661), .A2(P2_U3088), .ZN(n14205) );
  AOI22_X1 U12562 ( .A1(n14707), .A2(n10662), .B1(n14205), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n10663) );
  OAI211_X1 U12563 ( .C1(n10665), .C2(n11464), .A(n10664), .B(n10663), .ZN(
        P2_U3204) );
  INV_X1 U12564 ( .A(n10666), .ZN(n10673) );
  NAND3_X1 U12565 ( .A1(n14671), .A2(n14733), .A3(n10667), .ZN(n10668) );
  OAI21_X1 U12566 ( .B1(n14168), .B2(n14686), .A(n10668), .ZN(n10672) );
  AOI22_X1 U12567 ( .A1(n14911), .A2(n14733), .B1(n14731), .B2(n14913), .ZN(
        n10819) );
  INV_X1 U12568 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10669) );
  OAI22_X1 U12569 ( .A1(n14650), .A2(n10819), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10669), .ZN(n10671) );
  INV_X1 U12570 ( .A(n10998), .ZN(n16475) );
  OAI22_X1 U12571 ( .A1(n16472), .A2(n14683), .B1(n14705), .B2(n16475), .ZN(
        n10670) );
  AOI211_X1 U12572 ( .C1(n10673), .C2(n10672), .A(n10671), .B(n10670), .ZN(
        n10674) );
  OAI21_X1 U12573 ( .B1(n14686), .B2(n10723), .A(n10674), .ZN(P2_U3202) );
  XNOR2_X1 U12574 ( .A(n10830), .B(n11960), .ZN(n10677) );
  NOR2_X1 U12575 ( .A1(n10677), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10832) );
  AOI21_X1 U12576 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n10677), .A(n10832), 
        .ZN(n10686) );
  INV_X1 U12577 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10835) );
  MUX2_X1 U12578 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n10835), .S(n11960), .Z(
        n10680) );
  AOI21_X1 U12579 ( .B1(n11863), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10678), 
        .ZN(n10679) );
  NAND2_X1 U12580 ( .A1(n10679), .A2(n10680), .ZN(n10838) );
  OAI21_X1 U12581 ( .B1(n10680), .B2(n10679), .A(n10838), .ZN(n10684) );
  INV_X1 U12582 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n16288) );
  NAND2_X1 U12583 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n10682)
         );
  NAND2_X1 U12584 ( .A1(n15477), .A2(n11960), .ZN(n10681) );
  OAI211_X1 U12585 ( .C1(n15524), .C2(n16288), .A(n10682), .B(n10681), .ZN(
        n10683) );
  AOI21_X1 U12586 ( .B1(n10684), .B2(n15516), .A(n10683), .ZN(n10685) );
  OAI21_X1 U12587 ( .B1(n10686), .B2(n15398), .A(n10685), .ZN(P1_U3255) );
  INV_X1 U12588 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n10688) );
  NAND2_X1 U12589 ( .A1(n12618), .A2(n11644), .ZN(n10687) );
  OAI21_X1 U12590 ( .B1(P3_U3897), .B2(n10688), .A(n10687), .ZN(P3_U3502) );
  OAI21_X1 U12591 ( .B1(n10691), .B2(n10690), .A(n10689), .ZN(n11838) );
  XOR2_X1 U12592 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n11837), .Z(n10692) );
  XNOR2_X1 U12593 ( .A(n11838), .B(n10692), .ZN(n10706) );
  INV_X1 U12594 ( .A(n11837), .ZN(n10701) );
  INV_X1 U12595 ( .A(n10693), .ZN(n10695) );
  AOI21_X1 U12596 ( .B1(n10701), .B2(P2_REG1_REG_14__SCAN_IN), .A(n10695), 
        .ZN(n10694) );
  OAI21_X1 U12597 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n10701), .A(n10694), 
        .ZN(n10699) );
  NOR2_X1 U12598 ( .A1(n11837), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n10697) );
  NOR2_X1 U12599 ( .A1(n10700), .A2(n10695), .ZN(n10696) );
  AOI211_X1 U12600 ( .C1(n11837), .C2(P2_REG1_REG_14__SCAN_IN), .A(n10697), 
        .B(n10696), .ZN(n11825) );
  INV_X1 U12601 ( .A(n11825), .ZN(n10698) );
  OAI211_X1 U12602 ( .C1(n10700), .C2(n10699), .A(n10698), .B(n16148), .ZN(
        n10705) );
  NOR2_X1 U12603 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n12129), .ZN(n10703) );
  NOR2_X1 U12604 ( .A1(n16127), .A2(n10701), .ZN(n10702) );
  AOI211_X1 U12605 ( .C1(n16110), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n10703), 
        .B(n10702), .ZN(n10704) );
  OAI211_X1 U12606 ( .C1(n10706), .C2(n16114), .A(n10705), .B(n10704), .ZN(
        P2_U3228) );
  INV_X1 U12607 ( .A(n14205), .ZN(n10709) );
  OAI22_X1 U12608 ( .A1(n10709), .A2(n10708), .B1(n10707), .B2(n14650), .ZN(
        n10715) );
  AOI22_X1 U12609 ( .A1(n14671), .A2(n14735), .B1(n14707), .B2(n10710), .ZN(
        n10713) );
  INV_X1 U12610 ( .A(n10711), .ZN(n14203) );
  NOR3_X1 U12611 ( .A1(n10713), .A2(n14203), .A3(n10712), .ZN(n10714) );
  AOI211_X1 U12612 ( .C1(n10716), .C2(n14691), .A(n10715), .B(n10714), .ZN(
        n10717) );
  OAI21_X1 U12613 ( .B1(n14686), .B2(n10718), .A(n10717), .ZN(P2_U3209) );
  INV_X1 U12614 ( .A(n14650), .ZN(n14681) );
  OAI22_X1 U12615 ( .A1(n11350), .A2(n14953), .B1(n10997), .B2(n14951), .ZN(
        n11001) );
  AND2_X1 U12616 ( .A1(n14681), .A2(n11001), .ZN(n10720) );
  INV_X1 U12617 ( .A(n11802), .ZN(n11347) );
  OAI22_X1 U12618 ( .A1(n14683), .A2(n11799), .B1(n14705), .B2(n11347), .ZN(
        n10719) );
  AOI211_X1 U12619 ( .C1(P2_REG3_REG_5__SCAN_IN), .C2(P2_U3088), .A(n10720), 
        .B(n10719), .ZN(n10726) );
  OAI22_X1 U12620 ( .A1(n10997), .A2(n14694), .B1(n14686), .B2(n10721), .ZN(
        n10724) );
  NAND3_X1 U12621 ( .A1(n10724), .A2(n8045), .A3(n10723), .ZN(n10725) );
  OAI211_X1 U12622 ( .C1(n10727), .C2(n14686), .A(n10726), .B(n10725), .ZN(
        P2_U3199) );
  INV_X1 U12623 ( .A(n11032), .ZN(n11528) );
  NAND2_X1 U12624 ( .A1(n10636), .A2(n11528), .ZN(n12787) );
  AND2_X1 U12625 ( .A1(n11537), .A2(n12787), .ZN(n12926) );
  AND2_X1 U12626 ( .A1(n10728), .A2(n16580), .ZN(n10729) );
  NAND2_X1 U12627 ( .A1(n10743), .A2(n10729), .ZN(n10731) );
  OR2_X1 U12628 ( .A1(n10746), .A2(n10738), .ZN(n10730) );
  NAND2_X1 U12629 ( .A1(n10731), .A2(n10730), .ZN(n10733) );
  INV_X1 U12630 ( .A(n10746), .ZN(n11039) );
  NOR2_X1 U12631 ( .A1(n11165), .A2(n10929), .ZN(n12961) );
  NAND3_X1 U12632 ( .A1(n11039), .A2(n12961), .A3(n11037), .ZN(n13593) );
  INV_X1 U12633 ( .A(n10743), .ZN(n10735) );
  INV_X1 U12634 ( .A(n12920), .ZN(n11534) );
  NAND2_X1 U12635 ( .A1(n10735), .A2(n11534), .ZN(n10736) );
  NOR2_X1 U12636 ( .A1(n10929), .A2(n16580), .ZN(n11522) );
  AOI22_X1 U12637 ( .A1(n10734), .A2(n13566), .B1(n13596), .B2(n11032), .ZN(
        n10750) );
  AND2_X1 U12638 ( .A1(n11513), .A2(n10737), .ZN(n10741) );
  INV_X1 U12639 ( .A(n10738), .ZN(n10739) );
  NAND2_X1 U12640 ( .A1(n10746), .A2(n10739), .ZN(n10740) );
  OAI211_X1 U12641 ( .C1(n10743), .C2(n10742), .A(n10741), .B(n10740), .ZN(
        n10744) );
  NAND2_X1 U12642 ( .A1(n10744), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10748) );
  OR2_X1 U12643 ( .A1(n10926), .A2(P3_U3151), .ZN(n12965) );
  INV_X1 U12644 ( .A(n12965), .ZN(n10745) );
  AOI21_X1 U12645 ( .B1(n12961), .B2(n10746), .A(n10745), .ZN(n10747) );
  NAND2_X1 U12646 ( .A1(n13448), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11199) );
  NAND2_X1 U12647 ( .A1(n11199), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10749) );
  OAI211_X1 U12648 ( .C1(n12926), .C2(n13599), .A(n10750), .B(n10749), .ZN(
        P3_U3172) );
  INV_X1 U12649 ( .A(n10751), .ZN(n10753) );
  NAND2_X1 U12650 ( .A1(n10753), .A2(n10752), .ZN(n10763) );
  NAND2_X1 U12651 ( .A1(n10765), .A2(n10763), .ZN(n10761) );
  OR2_X1 U12652 ( .A1(n10878), .A2(n15223), .ZN(n10759) );
  NAND2_X1 U12653 ( .A1(n10754), .A2(n13289), .ZN(n10757) );
  AOI22_X1 U12654 ( .A1(n13155), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n13154), 
        .B2(n10755), .ZN(n10756) );
  NAND2_X1 U12655 ( .A1(n10757), .A2(n10756), .ZN(n11362) );
  NAND2_X1 U12656 ( .A1(n11362), .A2(n7432), .ZN(n10758) );
  AND2_X1 U12657 ( .A1(n10759), .A2(n10758), .ZN(n10762) );
  INV_X1 U12658 ( .A(n10762), .ZN(n10760) );
  AND2_X1 U12659 ( .A1(n10763), .A2(n10762), .ZN(n10764) );
  NAND2_X1 U12660 ( .A1(n10765), .A2(n10764), .ZN(n10782) );
  NAND2_X1 U12661 ( .A1(n10783), .A2(n10782), .ZN(n10768) );
  NAND2_X1 U12662 ( .A1(n11362), .A2(n15255), .ZN(n10766) );
  OAI21_X1 U12663 ( .B1(n10878), .B2(n7462), .A(n10766), .ZN(n10767) );
  XNOR2_X1 U12664 ( .A(n10767), .B(n15253), .ZN(n10781) );
  XNOR2_X1 U12665 ( .A(n10768), .B(n10781), .ZN(n10779) );
  NAND2_X1 U12666 ( .A1(n13170), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n10774) );
  OR2_X1 U12667 ( .A1(n13256), .A2(n10769), .ZN(n10773) );
  NAND2_X1 U12668 ( .A1(n10770), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10799) );
  OAI21_X1 U12669 ( .B1(n10770), .B2(P1_REG3_REG_5__SCAN_IN), .A(n10799), .ZN(
        n11185) );
  OR2_X1 U12670 ( .A1(n13282), .A2(n11185), .ZN(n10772) );
  OR2_X1 U12671 ( .A1(n13284), .A2(n10437), .ZN(n10771) );
  INV_X1 U12672 ( .A(n15380), .ZN(n11204) );
  OAI22_X1 U12673 ( .A1(n11204), .A2(n15362), .B1(n15359), .B2(n10876), .ZN(
        n10778) );
  NAND2_X1 U12674 ( .A1(n15365), .A2(n11362), .ZN(n10776) );
  OAI211_X1 U12675 ( .C1(n15360), .C2(n11367), .A(n10776), .B(n10775), .ZN(
        n10777) );
  AOI211_X1 U12676 ( .C1(n10779), .C2(n15332), .A(n10778), .B(n10777), .ZN(
        n10780) );
  INV_X1 U12677 ( .A(n10780), .ZN(P1_U3230) );
  NAND2_X1 U12678 ( .A1(n15380), .A2(n7432), .ZN(n10788) );
  NAND2_X1 U12679 ( .A1(n10784), .A2(n13289), .ZN(n10786) );
  AOI22_X1 U12680 ( .A1(n13155), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n13154), 
        .B2(n15431), .ZN(n10785) );
  NAND2_X1 U12681 ( .A1(n10786), .A2(n10785), .ZN(n13053) );
  NAND2_X1 U12682 ( .A1(n13053), .A2(n15255), .ZN(n10787) );
  NAND2_X1 U12683 ( .A1(n10788), .A2(n10787), .ZN(n10789) );
  XNOR2_X1 U12684 ( .A(n10789), .B(n15253), .ZN(n10792) );
  OR2_X1 U12685 ( .A1(n11204), .A2(n15223), .ZN(n10791) );
  NAND2_X1 U12686 ( .A1(n13053), .A2(n7432), .ZN(n10790) );
  NAND2_X1 U12687 ( .A1(n10791), .A2(n10790), .ZN(n10793) );
  INV_X1 U12688 ( .A(n10792), .ZN(n10795) );
  INV_X1 U12689 ( .A(n10793), .ZN(n10794) );
  NAND2_X1 U12690 ( .A1(n10795), .A2(n10794), .ZN(n10891) );
  NAND2_X1 U12691 ( .A1(n7568), .A2(n10891), .ZN(n10796) );
  XNOR2_X1 U12692 ( .A(n10890), .B(n10796), .ZN(n10809) );
  NAND2_X1 U12693 ( .A1(n13277), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10805) );
  OR2_X1 U12694 ( .A1(n13284), .A2(n16496), .ZN(n10804) );
  AND2_X1 U12695 ( .A1(n10799), .A2(n10798), .ZN(n10800) );
  OR2_X1 U12696 ( .A1(n10800), .A2(n10902), .ZN(n11215) );
  OR2_X1 U12697 ( .A1(n13282), .A2(n11215), .ZN(n10803) );
  INV_X1 U12698 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10801) );
  OR2_X1 U12699 ( .A1(n13279), .A2(n10801), .ZN(n10802) );
  NAND4_X1 U12700 ( .A1(n10805), .A2(n10804), .A3(n10803), .A4(n10802), .ZN(
        n15379) );
  INV_X1 U12701 ( .A(n15379), .ZN(n11065) );
  OAI22_X1 U12702 ( .A1(n10878), .A2(n15359), .B1(n15362), .B2(n11065), .ZN(
        n10808) );
  NAND2_X1 U12703 ( .A1(n15365), .A2(n13053), .ZN(n10806) );
  NAND2_X1 U12704 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n15424) );
  OAI211_X1 U12705 ( .C1(n15360), .C2(n11185), .A(n10806), .B(n15424), .ZN(
        n10807) );
  AOI211_X1 U12706 ( .C1(n10809), .C2(n15332), .A(n10808), .B(n10807), .ZN(
        n10810) );
  INV_X1 U12707 ( .A(n10810), .ZN(P1_U3227) );
  NAND2_X1 U12708 ( .A1(n10812), .A2(n10811), .ZN(n10814) );
  INV_X1 U12709 ( .A(n14733), .ZN(n10817) );
  NAND2_X1 U12710 ( .A1(n11990), .A2(n10817), .ZN(n10813) );
  NAND2_X1 U12711 ( .A1(n10814), .A2(n10813), .ZN(n10991) );
  INV_X1 U12712 ( .A(n10995), .ZN(n10990) );
  XNOR2_X1 U12713 ( .A(n10991), .B(n10990), .ZN(n16478) );
  INV_X1 U12714 ( .A(n16478), .ZN(n10825) );
  NAND2_X1 U12715 ( .A1(n14170), .A2(n10817), .ZN(n10818) );
  XNOR2_X1 U12716 ( .A(n10996), .B(n10990), .ZN(n10820) );
  OAI21_X1 U12717 ( .B1(n10820), .B2(n14949), .A(n10819), .ZN(n10821) );
  AOI21_X1 U12718 ( .B1(n16507), .B2(n16478), .A(n10821), .ZN(n16481) );
  OR2_X1 U12719 ( .A1(n10823), .A2(n10998), .ZN(n10987) );
  INV_X1 U12720 ( .A(n10987), .ZN(n10822) );
  AOI211_X1 U12721 ( .C1(n10998), .C2(n10823), .A(n14986), .B(n10822), .ZN(
        n16477) );
  AOI21_X1 U12722 ( .B1(n15079), .B2(n10998), .A(n16477), .ZN(n10824) );
  OAI211_X1 U12723 ( .C1(n10450), .C2(n10825), .A(n16481), .B(n10824), .ZN(
        n15084) );
  NAND2_X1 U12724 ( .A1(n15084), .A2(n15102), .ZN(n10826) );
  OAI21_X1 U12725 ( .B1(n15102), .B2(n8640), .A(n10826), .ZN(P2_U3442) );
  INV_X1 U12726 ( .A(n10827), .ZN(n10828) );
  OAI222_X1 U12727 ( .A1(n14150), .A2(n10829), .B1(n14154), .B2(n10828), .C1(
        n13668), .C2(P3_U3151), .ZN(P3_U3278) );
  INV_X1 U12728 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11973) );
  XNOR2_X1 U12729 ( .A(n11445), .B(n11973), .ZN(n10834) );
  NOR2_X1 U12730 ( .A1(n10830), .A2(n11960), .ZN(n10831) );
  OR2_X1 U12731 ( .A1(n10832), .A2(n10831), .ZN(n10833) );
  NOR3_X1 U12732 ( .A1(n10832), .A2(n10831), .A3(n10834), .ZN(n11452) );
  AOI211_X1 U12733 ( .C1(n10834), .C2(n10833), .A(n15398), .B(n11452), .ZN(
        n10844) );
  NAND2_X1 U12734 ( .A1(n10836), .A2(n10835), .ZN(n10837) );
  AND2_X1 U12735 ( .A1(n10838), .A2(n10837), .ZN(n10840) );
  XNOR2_X1 U12736 ( .A(n11445), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n10839) );
  NAND3_X1 U12737 ( .A1(n10838), .A2(n10839), .A3(n10837), .ZN(n11449) );
  OAI211_X1 U12738 ( .C1(n10840), .C2(n10839), .A(n15516), .B(n11449), .ZN(
        n10842) );
  AND2_X1 U12739 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n12365) );
  AOI21_X1 U12740 ( .B1(n16162), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n12365), 
        .ZN(n10841) );
  OAI211_X1 U12741 ( .C1(n15511), .C2(n11445), .A(n10842), .B(n10841), .ZN(
        n10843) );
  OR2_X1 U12742 ( .A1(n10844), .A2(n10843), .ZN(P1_U3256) );
  OAI222_X1 U12743 ( .A1(P3_U3151), .A2(n13680), .B1(n14150), .B2(n14425), 
        .C1(n14154), .C2(n10845), .ZN(P3_U3277) );
  NAND2_X1 U12744 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n14784) );
  OAI21_X1 U12745 ( .B1(n14683), .B2(n16510), .A(n14784), .ZN(n10847) );
  INV_X1 U12746 ( .A(n11548), .ZN(n16516) );
  OAI22_X1 U12747 ( .A1(n11464), .A2(n11551), .B1(n16516), .B2(n14705), .ZN(
        n10846) );
  AOI211_X1 U12748 ( .C1(n14701), .C2(n14730), .A(n10847), .B(n10846), .ZN(
        n10854) );
  NAND3_X1 U12749 ( .A1(n14671), .A2(n14730), .A3(n10848), .ZN(n10849) );
  OAI21_X1 U12750 ( .B1(n11045), .B2(n14686), .A(n10849), .ZN(n10852) );
  INV_X1 U12751 ( .A(n10850), .ZN(n10851) );
  NAND2_X1 U12752 ( .A1(n10852), .A2(n10851), .ZN(n10853) );
  OAI211_X1 U12753 ( .C1(n10855), .C2(n14686), .A(n10854), .B(n10853), .ZN(
        P2_U3185) );
  OR2_X1 U12754 ( .A1(n10856), .A2(P1_U3086), .ZN(n13366) );
  NAND3_X1 U12755 ( .A1(n10859), .A2(n10858), .A3(n10857), .ZN(n10860) );
  NOR2_X1 U12756 ( .A1(n13366), .A2(n10860), .ZN(n11054) );
  INV_X1 U12757 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10888) );
  NAND2_X1 U12758 ( .A1(n15384), .A2(n13025), .ZN(n10861) );
  NAND2_X1 U12759 ( .A1(n16434), .A2(n15383), .ZN(n13022) );
  NAND2_X1 U12760 ( .A1(n11137), .A2(n10875), .ZN(n10864) );
  NAND2_X1 U12761 ( .A1(n7856), .A2(n16434), .ZN(n10863) );
  NAND2_X1 U12762 ( .A1(n10864), .A2(n10863), .ZN(n11172) );
  INV_X1 U12763 ( .A(n10876), .ZN(n15382) );
  INV_X1 U12764 ( .A(n13312), .ZN(n10865) );
  NAND2_X1 U12765 ( .A1(n11172), .A2(n10865), .ZN(n10867) );
  NAND2_X1 U12766 ( .A1(n16452), .A2(n10876), .ZN(n10866) );
  AND2_X1 U12767 ( .A1(n16463), .A2(n10878), .ZN(n10869) );
  OR2_X1 U12768 ( .A1(n16463), .A2(n10878), .ZN(n10868) );
  INV_X1 U12769 ( .A(n13311), .ZN(n11063) );
  XNOR2_X1 U12770 ( .A(n11064), .B(n11063), .ZN(n11190) );
  OR2_X1 U12771 ( .A1(n10870), .A2(n13028), .ZN(n10871) );
  NAND2_X1 U12772 ( .A1(n11136), .A2(n15519), .ZN(n16454) );
  INV_X1 U12773 ( .A(n13310), .ZN(n10873) );
  OR2_X1 U12774 ( .A1(n15384), .A2(n7601), .ZN(n10874) );
  NAND2_X1 U12775 ( .A1(n11125), .A2(n10874), .ZN(n11139) );
  INV_X1 U12776 ( .A(n10875), .ZN(n13313) );
  NAND2_X1 U12777 ( .A1(n11139), .A2(n13313), .ZN(n11138) );
  NAND2_X1 U12778 ( .A1(n11138), .A2(n13021), .ZN(n11180) );
  NAND2_X1 U12779 ( .A1(n16452), .A2(n15382), .ZN(n13043) );
  NAND2_X1 U12780 ( .A1(n11180), .A2(n13043), .ZN(n10877) );
  NAND2_X1 U12781 ( .A1(n10876), .A2(n11173), .ZN(n13042) );
  AND2_X1 U12782 ( .A1(n10878), .A2(n11362), .ZN(n13048) );
  INV_X1 U12783 ( .A(n10878), .ZN(n15381) );
  NAND2_X1 U12784 ( .A1(n16463), .A2(n15381), .ZN(n13050) );
  XNOR2_X1 U12785 ( .A(n11055), .B(n11063), .ZN(n10881) );
  OR2_X1 U12786 ( .A1(n12983), .A2(n15519), .ZN(n10880) );
  NAND2_X1 U12787 ( .A1(n12984), .A2(n12998), .ZN(n10879) );
  NAND2_X1 U12788 ( .A1(n10881), .A2(n16458), .ZN(n10883) );
  AOI22_X1 U12789 ( .A1(n15381), .A2(n15787), .B1(n15789), .B2(n15379), .ZN(
        n10882) );
  OAI211_X1 U12790 ( .C1(n11190), .C2(n16454), .A(n10883), .B(n10882), .ZN(
        n11183) );
  INV_X1 U12791 ( .A(n11183), .ZN(n10886) );
  NAND2_X1 U12792 ( .A1(n16434), .A2(n11142), .ZN(n11174) );
  INV_X1 U12793 ( .A(n11366), .ZN(n10884) );
  INV_X1 U12794 ( .A(n13053), .ZN(n13054) );
  AOI211_X1 U12795 ( .C1(n13053), .C2(n10884), .A(n15915), .B(n11211), .ZN(
        n11187) );
  AOI21_X1 U12796 ( .B1(n16490), .B2(n13053), .A(n11187), .ZN(n10885) );
  OAI211_X1 U12797 ( .C1(n11190), .C2(n16493), .A(n10886), .B(n10885), .ZN(
        n15945) );
  NAND2_X1 U12798 ( .A1(n15945), .A2(n16570), .ZN(n10887) );
  OAI21_X1 U12799 ( .B1(n16570), .B2(n10888), .A(n10887), .ZN(P1_U3474) );
  INV_X1 U12800 ( .A(n13109), .ZN(n11011) );
  INV_X1 U12801 ( .A(n11836), .ZN(n16086) );
  OAI222_X1 U12802 ( .A1(n15131), .A2(n11011), .B1(n16086), .B2(P2_U3088), 
        .C1(n10889), .C2(n15133), .ZN(P2_U3311) );
  OR2_X1 U12803 ( .A1(n10892), .A2(n12973), .ZN(n10895) );
  AOI22_X1 U12804 ( .A1(n13155), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n13154), 
        .B2(n10893), .ZN(n10894) );
  NAND2_X1 U12805 ( .A1(n10895), .A2(n10894), .ZN(n16489) );
  NAND2_X1 U12806 ( .A1(n16489), .A2(n15255), .ZN(n10897) );
  NAND2_X1 U12807 ( .A1(n15379), .A2(n7432), .ZN(n10896) );
  NAND2_X1 U12808 ( .A1(n10897), .A2(n10896), .ZN(n10898) );
  XNOR2_X1 U12809 ( .A(n10898), .B(n15221), .ZN(n11105) );
  NAND2_X1 U12810 ( .A1(n16489), .A2(n7432), .ZN(n10900) );
  OR2_X1 U12811 ( .A1(n11065), .A2(n15223), .ZN(n10899) );
  AND2_X1 U12812 ( .A1(n10900), .A2(n10899), .ZN(n11103) );
  INV_X1 U12813 ( .A(n11103), .ZN(n11106) );
  XNOR2_X1 U12814 ( .A(n11105), .B(n11106), .ZN(n10901) );
  XNOR2_X1 U12815 ( .A(n11104), .B(n10901), .ZN(n10912) );
  NAND2_X1 U12816 ( .A1(n13170), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n10907) );
  OR2_X1 U12817 ( .A1(n13256), .A2(n11331), .ZN(n10906) );
  NAND2_X1 U12818 ( .A1(n10902), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11071) );
  OR2_X1 U12819 ( .A1(n10902), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10903) );
  NAND2_X1 U12820 ( .A1(n11071), .A2(n10903), .ZN(n11333) );
  OR2_X1 U12821 ( .A1(n13282), .A2(n11333), .ZN(n10905) );
  OR2_X1 U12822 ( .A1(n13284), .A2(n11082), .ZN(n10904) );
  NAND4_X1 U12823 ( .A1(n10907), .A2(n10906), .A3(n10905), .A4(n10904), .ZN(
        n15378) );
  INV_X1 U12824 ( .A(n15378), .ZN(n11566) );
  OAI22_X1 U12825 ( .A1(n11566), .A2(n15362), .B1(n15359), .B2(n11204), .ZN(
        n10911) );
  NAND2_X1 U12826 ( .A1(n15365), .A2(n16489), .ZN(n10909) );
  OAI211_X1 U12827 ( .C1(n15360), .C2(n11215), .A(n10909), .B(n10908), .ZN(
        n10910) );
  AOI211_X1 U12828 ( .C1(n10912), .C2(n15332), .A(n10911), .B(n10910), .ZN(
        n10913) );
  INV_X1 U12829 ( .A(n10913), .ZN(P1_U3239) );
  MUX2_X1 U12830 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n13671), .Z(n10915) );
  XOR2_X1 U12831 ( .A(n14155), .B(n10915), .Z(n11013) );
  INV_X1 U12832 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11525) );
  MUX2_X1 U12833 ( .A(n11525), .B(n9586), .S(n13671), .Z(n11147) );
  NAND2_X1 U12834 ( .A1(n11147), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11146) );
  INV_X1 U12835 ( .A(n14155), .ZN(n10914) );
  OAI22_X1 U12836 ( .A1(n11013), .A2(n11146), .B1(n10915), .B2(n10914), .ZN(
        n11086) );
  MUX2_X1 U12837 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n13671), .Z(n10916) );
  XOR2_X1 U12838 ( .A(n7619), .B(n10916), .Z(n11087) );
  INV_X1 U12839 ( .A(n7619), .ZN(n10918) );
  INV_X1 U12840 ( .A(n10916), .ZN(n10917) );
  AOI22_X1 U12841 ( .A1(n11086), .A2(n11087), .B1(n10918), .B2(n10917), .ZN(
        n11267) );
  MUX2_X1 U12842 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n7429), .Z(n10919) );
  XOR2_X1 U12843 ( .A(n11277), .B(n10919), .Z(n11268) );
  INV_X1 U12844 ( .A(n11277), .ZN(n10949) );
  OAI22_X1 U12845 ( .A1(n11267), .A2(n11268), .B1(n10919), .B2(n10949), .ZN(
        n11249) );
  MUX2_X1 U12846 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n7429), .Z(n10920) );
  XNOR2_X1 U12847 ( .A(n10920), .B(n10953), .ZN(n11248) );
  INV_X1 U12848 ( .A(n10920), .ZN(n10921) );
  MUX2_X1 U12849 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n7429), .Z(n10922) );
  XNOR2_X1 U12850 ( .A(n10922), .B(n10955), .ZN(n10973) );
  MUX2_X1 U12851 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n7429), .Z(n10923) );
  NOR2_X1 U12852 ( .A1(n10923), .A2(n11226), .ZN(n11222) );
  INV_X1 U12853 ( .A(n11222), .ZN(n10924) );
  NAND2_X1 U12854 ( .A1(n10923), .A2(n11226), .ZN(n11221) );
  NAND2_X1 U12855 ( .A1(n10924), .A2(n11221), .ZN(n10925) );
  XNOR2_X1 U12856 ( .A(n11223), .B(n10925), .ZN(n10971) );
  NAND2_X1 U12857 ( .A1(P3_U3897), .A2(n12732), .ZN(n16376) );
  NAND2_X1 U12858 ( .A1(n12910), .A2(n10926), .ZN(n10927) );
  NAND2_X1 U12859 ( .A1(n10928), .A2(n10927), .ZN(n10962) );
  AND2_X1 U12860 ( .A1(n10929), .A2(n12965), .ZN(n10961) );
  NOR2_X1 U12861 ( .A1(n10962), .A2(n10961), .ZN(n10960) );
  INV_X1 U12862 ( .A(n10930), .ZN(n10931) );
  NAND2_X1 U12863 ( .A1(n10960), .A2(n10931), .ZN(n16382) );
  MUX2_X1 U12864 ( .A(P3_REG2_REG_2__SCAN_IN), .B(n10932), .S(n11097), .Z(
        n11090) );
  AND2_X1 U12865 ( .A1(n9615), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10934) );
  NAND2_X1 U12866 ( .A1(n11152), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10933) );
  OAI22_X1 U12867 ( .A1(n10934), .A2(n14155), .B1(n9615), .B2(n10933), .ZN(
        n11014) );
  NAND2_X1 U12868 ( .A1(n11014), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n10936) );
  INV_X1 U12869 ( .A(n10934), .ZN(n10935) );
  NAND2_X1 U12870 ( .A1(n10936), .A2(n10935), .ZN(n11089) );
  NAND2_X1 U12871 ( .A1(n7619), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10937) );
  NAND2_X1 U12872 ( .A1(n11088), .A2(n10937), .ZN(n10938) );
  NAND2_X1 U12873 ( .A1(n11269), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n10940) );
  NAND2_X1 U12874 ( .A1(n10938), .A2(n10949), .ZN(n10939) );
  NAND2_X1 U12875 ( .A1(n10940), .A2(n10939), .ZN(n11252) );
  MUX2_X1 U12876 ( .A(n10941), .B(P3_REG2_REG_4__SCAN_IN), .S(n10953), .Z(
        n11253) );
  NAND2_X1 U12877 ( .A1(n11252), .A2(n11253), .ZN(n11251) );
  OAI21_X1 U12878 ( .B1(n10953), .B2(n10941), .A(n11251), .ZN(n10942) );
  XNOR2_X1 U12879 ( .A(n10942), .B(n10955), .ZN(n10974) );
  INV_X1 U12880 ( .A(n10942), .ZN(n10943) );
  INV_X1 U12881 ( .A(n10955), .ZN(n10978) );
  XNOR2_X1 U12882 ( .A(n11230), .B(P3_REG2_REG_6__SCAN_IN), .ZN(n11227) );
  XNOR2_X1 U12883 ( .A(n11228), .B(n11227), .ZN(n10969) );
  INV_X1 U12884 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n16428) );
  NAND2_X1 U12885 ( .A1(n11152), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10945) );
  NAND2_X1 U12886 ( .A1(n14155), .A2(n10945), .ZN(n10946) );
  NAND2_X1 U12887 ( .A1(n9615), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10947) );
  NAND2_X1 U12888 ( .A1(n10946), .A2(n10947), .ZN(n11016) );
  INV_X1 U12889 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n16405) );
  OR2_X1 U12890 ( .A1(n11016), .A2(n16405), .ZN(n11018) );
  NAND2_X1 U12891 ( .A1(n11018), .A2(n10947), .ZN(n11092) );
  NAND2_X1 U12892 ( .A1(n7619), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10948) );
  NAND2_X1 U12893 ( .A1(n10950), .A2(n10949), .ZN(n11257) );
  OAI21_X1 U12894 ( .B1(n10950), .B2(n10949), .A(n11257), .ZN(n11270) );
  INV_X1 U12895 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n16448) );
  OR2_X1 U12896 ( .A1(n11270), .A2(n16448), .ZN(n11272) );
  NAND2_X1 U12897 ( .A1(n11272), .A2(n11257), .ZN(n10952) );
  INV_X1 U12898 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10951) );
  MUX2_X1 U12899 ( .A(n10951), .B(P3_REG1_REG_4__SCAN_IN), .S(n10953), .Z(
        n11256) );
  NAND2_X1 U12900 ( .A1(n10952), .A2(n11256), .ZN(n11260) );
  INV_X1 U12901 ( .A(n10953), .ZN(n11266) );
  NAND2_X1 U12902 ( .A1(n11266), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10954) );
  NAND2_X1 U12903 ( .A1(n11260), .A2(n10954), .ZN(n10956) );
  INV_X1 U12904 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n16486) );
  XNOR2_X1 U12905 ( .A(n11230), .B(P3_REG1_REG_6__SCAN_IN), .ZN(n10957) );
  INV_X1 U12906 ( .A(n10957), .ZN(n10958) );
  AND2_X1 U12907 ( .A1(n11232), .A2(n10959), .ZN(n10967) );
  NAND2_X1 U12908 ( .A1(n10960), .A2(n7429), .ZN(n16374) );
  MUX2_X1 U12909 ( .A(n10960), .B(P3_U3897), .S(n12960), .Z(n13707) );
  NAND2_X1 U12910 ( .A1(n13707), .A2(n11230), .ZN(n10966) );
  INV_X1 U12911 ( .A(n10961), .ZN(n10963) );
  INV_X1 U12912 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10964) );
  NOR2_X1 U12913 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10964), .ZN(n12162) );
  AOI21_X1 U12914 ( .B1(n16036), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n12162), .ZN(
        n10965) );
  OAI211_X1 U12915 ( .C1(n10967), .C2(n16374), .A(n10966), .B(n10965), .ZN(
        n10968) );
  AOI21_X1 U12916 ( .B1(n13712), .B2(n10969), .A(n10968), .ZN(n10970) );
  OAI21_X1 U12917 ( .B1(n10971), .B2(n16376), .A(n10970), .ZN(P3_U3188) );
  XOR2_X1 U12918 ( .A(n10972), .B(n10973), .Z(n10986) );
  XOR2_X1 U12919 ( .A(n10974), .B(P3_REG2_REG_5__SCAN_IN), .Z(n10984) );
  NAND2_X1 U12920 ( .A1(n10975), .A2(n16486), .ZN(n10976) );
  AND2_X1 U12921 ( .A1(n10977), .A2(n10976), .ZN(n10982) );
  NAND2_X1 U12922 ( .A1(n13707), .A2(n10978), .ZN(n10981) );
  INV_X1 U12923 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10979) );
  NOR2_X1 U12924 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10979), .ZN(n11714) );
  AOI21_X1 U12925 ( .B1(n16036), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11714), .ZN(
        n10980) );
  OAI211_X1 U12926 ( .C1(n10982), .C2(n16374), .A(n10981), .B(n10980), .ZN(
        n10983) );
  AOI21_X1 U12927 ( .B1(n13712), .B2(n10984), .A(n10983), .ZN(n10985) );
  OAI21_X1 U12928 ( .B1(n10986), .B2(n16376), .A(n10985), .ZN(P3_U3187) );
  NAND2_X1 U12929 ( .A1(n10987), .A2(n11802), .ZN(n10988) );
  NAND2_X1 U12930 ( .A1(n10988), .A2(n14930), .ZN(n10989) );
  NOR2_X1 U12931 ( .A1(n11927), .A2(n10989), .ZN(n11798) );
  NAND2_X1 U12932 ( .A1(n10991), .A2(n10990), .ZN(n10993) );
  OR2_X1 U12933 ( .A1(n14732), .A2(n10998), .ZN(n10992) );
  NAND2_X1 U12934 ( .A1(n10993), .A2(n10992), .ZN(n11341) );
  XNOR2_X1 U12935 ( .A(n11341), .B(n11000), .ZN(n11805) );
  NOR2_X1 U12936 ( .A1(n11805), .A2(n15082), .ZN(n10994) );
  AOI211_X1 U12937 ( .C1(n15079), .C2(n11802), .A(n11798), .B(n10994), .ZN(
        n11003) );
  NAND2_X1 U12938 ( .A1(n10998), .A2(n10997), .ZN(n10999) );
  XNOR2_X1 U12939 ( .A(n11346), .B(n11000), .ZN(n11002) );
  AOI21_X1 U12940 ( .B1(n11002), .B2(n14981), .A(n11001), .ZN(n11797) );
  NAND2_X1 U12941 ( .A1(n11003), .A2(n11797), .ZN(n11005) );
  NAND2_X1 U12942 ( .A1(n11005), .A2(n7433), .ZN(n11004) );
  OAI21_X1 U12943 ( .B1(n7433), .B2(n10289), .A(n11004), .ZN(P2_U3504) );
  NAND2_X1 U12944 ( .A1(n11005), .A2(n15102), .ZN(n11006) );
  OAI21_X1 U12945 ( .B1(n15102), .B2(n8661), .A(n11006), .ZN(P2_U3445) );
  INV_X1 U12946 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n11008) );
  NAND2_X1 U12947 ( .A1(n13794), .A2(n11644), .ZN(n11007) );
  OAI21_X1 U12948 ( .B1(P3_U3897), .B2(n11008), .A(n11007), .ZN(P3_U3514) );
  NAND2_X1 U12949 ( .A1(n11009), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11010) );
  XNOR2_X1 U12950 ( .A(n11010), .B(P1_IR_REG_16__SCAN_IN), .ZN(n13110) );
  INV_X1 U12951 ( .A(n13110), .ZN(n12340) );
  OAI222_X1 U12952 ( .A1(n15987), .A2(n11012), .B1(n15990), .B2(n11011), .C1(
        P1_U3086), .C2(n12340), .ZN(P1_U3339) );
  XOR2_X1 U12953 ( .A(n11013), .B(n11146), .Z(n11024) );
  XNOR2_X1 U12954 ( .A(n11014), .B(n11536), .ZN(n11015) );
  NOR2_X1 U12955 ( .A1(n16382), .A2(n11015), .ZN(n11022) );
  NAND2_X1 U12956 ( .A1(n11016), .A2(n16405), .ZN(n11017) );
  AND2_X1 U12957 ( .A1(n11018), .A2(n11017), .ZN(n11020) );
  AOI22_X1 U12958 ( .A1(n16036), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n11019) );
  OAI21_X1 U12959 ( .B1(n11020), .B2(n16374), .A(n11019), .ZN(n11021) );
  AOI211_X1 U12960 ( .C1(n13707), .C2(n14155), .A(n11022), .B(n11021), .ZN(
        n11023) );
  OAI21_X1 U12961 ( .B1(n16376), .B2(n11024), .A(n11023), .ZN(P3_U3183) );
  NAND2_X1 U12962 ( .A1(n11025), .A2(n11281), .ZN(n11030) );
  INV_X1 U12963 ( .A(n12953), .ZN(n11027) );
  NAND3_X1 U12964 ( .A1(n11028), .A2(n11027), .A3(n11026), .ZN(n11029) );
  OAI21_X1 U12965 ( .B1(n13425), .B2(n11032), .A(n11031), .ZN(n11036) );
  XNOR2_X1 U12966 ( .A(n11033), .B(n11499), .ZN(n11034) );
  OAI21_X1 U12967 ( .B1(n11654), .B2(n11034), .A(n11191), .ZN(n11035) );
  AOI21_X1 U12968 ( .B1(n11036), .B2(n11035), .A(n11193), .ZN(n11044) );
  INV_X1 U12969 ( .A(n12961), .ZN(n11038) );
  NOR2_X1 U12970 ( .A1(n11038), .A2(n11037), .ZN(n11040) );
  INV_X1 U12971 ( .A(n13568), .ZN(n13589) );
  AOI22_X1 U12972 ( .A1(n13566), .A2(n13483), .B1(n10636), .B2(n13589), .ZN(
        n11041) );
  OAI21_X1 U12973 ( .B1(n11529), .B2(n13582), .A(n11041), .ZN(n11042) );
  AOI21_X1 U12974 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(n11199), .A(n11042), .ZN(
        n11043) );
  OAI21_X1 U12975 ( .B1(n11044), .B2(n13599), .A(n11043), .ZN(P3_U3162) );
  INV_X1 U12976 ( .A(n11045), .ZN(n11046) );
  AOI211_X1 U12977 ( .C1(n11048), .C2(n11047), .A(n14686), .B(n11046), .ZN(
        n11052) );
  INV_X1 U12978 ( .A(n14701), .ZN(n11465) );
  INV_X1 U12979 ( .A(n14731), .ZN(n11344) );
  INV_X1 U12980 ( .A(n11934), .ZN(n16499) );
  OAI22_X1 U12981 ( .A1(n11465), .A2(n11344), .B1(n16499), .B2(n14705), .ZN(
        n11051) );
  NAND2_X1 U12982 ( .A1(n14702), .A2(n14729), .ZN(n11049) );
  NAND2_X1 U12983 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n14770) );
  OAI211_X1 U12984 ( .C1(n14683), .C2(n11930), .A(n11049), .B(n14770), .ZN(
        n11050) );
  OR3_X1 U12985 ( .A1(n11052), .A2(n11051), .A3(n11050), .ZN(P2_U3211) );
  INV_X1 U12986 ( .A(n11053), .ZN(n11118) );
  NAND2_X1 U12987 ( .A1(n13054), .A2(n15380), .ZN(n11056) );
  NAND2_X1 U12988 ( .A1(n11057), .A2(n11056), .ZN(n11205) );
  XNOR2_X1 U12989 ( .A(n16489), .B(n15379), .ZN(n13059) );
  NAND2_X1 U12990 ( .A1(n11205), .A2(n13059), .ZN(n11059) );
  INV_X1 U12991 ( .A(n16489), .ZN(n11216) );
  NAND2_X1 U12992 ( .A1(n11216), .A2(n15379), .ZN(n11058) );
  NAND2_X1 U12993 ( .A1(n11060), .A2(n13289), .ZN(n11062) );
  AOI22_X1 U12994 ( .A1(n13155), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n13154), 
        .B2(n15443), .ZN(n11061) );
  NAND2_X1 U12995 ( .A1(n11062), .A2(n11061), .ZN(n13065) );
  XNOR2_X1 U12996 ( .A(n13065), .B(n15378), .ZN(n13318) );
  XNOR2_X1 U12997 ( .A(n11568), .B(n13318), .ZN(n11340) );
  INV_X1 U12998 ( .A(n13059), .ZN(n13315) );
  NAND2_X1 U12999 ( .A1(n11216), .A2(n11065), .ZN(n11066) );
  NAND2_X1 U13000 ( .A1(n11202), .A2(n11066), .ZN(n11068) );
  INV_X1 U13001 ( .A(n13318), .ZN(n11067) );
  OAI21_X1 U13002 ( .B1(n11068), .B2(n11067), .A(n11562), .ZN(n11337) );
  INV_X1 U13003 ( .A(n13065), .ZN(n11329) );
  NAND2_X1 U13004 ( .A1(n13170), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n11076) );
  OR2_X1 U13005 ( .A1(n13256), .A2(n11069), .ZN(n11075) );
  OR2_X1 U13006 ( .A1(n13284), .A2(n11581), .ZN(n11074) );
  NAND2_X1 U13007 ( .A1(n11071), .A2(n11070), .ZN(n11072) );
  NAND2_X1 U13008 ( .A1(n11305), .A2(n11072), .ZN(n16523) );
  OR2_X1 U13009 ( .A1(n13282), .A2(n16523), .ZN(n11073) );
  NAND4_X1 U13010 ( .A1(n11076), .A2(n11075), .A3(n11074), .A4(n11073), .ZN(
        n15377) );
  NAND2_X1 U13011 ( .A1(n15789), .A2(n15377), .ZN(n11078) );
  NAND2_X1 U13012 ( .A1(n15787), .A2(n15379), .ZN(n11077) );
  AND2_X1 U13013 ( .A1(n11078), .A2(n11077), .ZN(n11330) );
  OAI21_X1 U13014 ( .B1(n11329), .B2(n16556), .A(n11330), .ZN(n11079) );
  OR2_X1 U13015 ( .A1(n11212), .A2(n13065), .ZN(n11572) );
  AOI211_X1 U13016 ( .C1(n13065), .C2(n11212), .A(n15915), .B(n7599), .ZN(
        n11336) );
  AOI211_X1 U13017 ( .C1(n11337), .C2(n16564), .A(n11079), .B(n11336), .ZN(
        n11080) );
  OAI21_X1 U13018 ( .B1(n16558), .B2(n11340), .A(n11080), .ZN(n11083) );
  NAND2_X1 U13019 ( .A1(n11083), .A2(n16469), .ZN(n11081) );
  OAI21_X1 U13020 ( .B1(n16469), .B2(n11082), .A(n11081), .ZN(P1_U3535) );
  INV_X1 U13021 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n11085) );
  NAND2_X1 U13022 ( .A1(n11083), .A2(n16570), .ZN(n11084) );
  OAI21_X1 U13023 ( .B1(n16570), .B2(n11085), .A(n11084), .ZN(P1_U3480) );
  XOR2_X1 U13024 ( .A(n11086), .B(n11087), .Z(n11102) );
  OAI21_X1 U13025 ( .B1(n11090), .B2(n11089), .A(n11088), .ZN(n11100) );
  OAI21_X1 U13026 ( .B1(n11093), .B2(n11092), .A(n11091), .ZN(n11094) );
  INV_X1 U13027 ( .A(n11094), .ZN(n11096) );
  AOI22_X1 U13028 ( .A1(n16036), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n11095) );
  OAI21_X1 U13029 ( .B1(n11096), .B2(n16374), .A(n11095), .ZN(n11099) );
  NOR2_X1 U13030 ( .A1(n16367), .A2(n7619), .ZN(n11098) );
  AOI211_X1 U13031 ( .C1(n13712), .C2(n11100), .A(n11099), .B(n11098), .ZN(
        n11101) );
  OAI21_X1 U13032 ( .B1(n11102), .B2(n16376), .A(n11101), .ZN(P3_U3184) );
  INV_X1 U13033 ( .A(n11105), .ZN(n11107) );
  NAND2_X1 U13034 ( .A1(n11107), .A2(n11106), .ZN(n11108) );
  NAND2_X1 U13035 ( .A1(n13065), .A2(n15255), .ZN(n11111) );
  NAND2_X1 U13036 ( .A1(n15378), .A2(n7432), .ZN(n11110) );
  NAND2_X1 U13037 ( .A1(n11111), .A2(n11110), .ZN(n11112) );
  XNOR2_X1 U13038 ( .A(n11112), .B(n15253), .ZN(n11286) );
  NOR2_X1 U13039 ( .A1(n11566), .A2(n15223), .ZN(n11113) );
  AOI21_X1 U13040 ( .B1(n13065), .B2(n7432), .A(n11113), .ZN(n11287) );
  XNOR2_X1 U13041 ( .A(n11286), .B(n11287), .ZN(n11284) );
  XNOR2_X1 U13042 ( .A(n11285), .B(n11284), .ZN(n11117) );
  NAND2_X1 U13043 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n15440) );
  OAI21_X1 U13044 ( .B1(n15264), .B2(n11330), .A(n15440), .ZN(n11115) );
  NOR2_X1 U13045 ( .A1(n15360), .A2(n11333), .ZN(n11114) );
  AOI211_X1 U13046 ( .C1(n13065), .C2(n15365), .A(n11115), .B(n11114), .ZN(
        n11116) );
  OAI21_X1 U13047 ( .B1(n11117), .B2(n15367), .A(n11116), .ZN(P1_U3213) );
  INV_X1 U13048 ( .A(n13366), .ZN(n11121) );
  NOR2_X1 U13049 ( .A1(n11119), .A2(n11118), .ZN(n11120) );
  NAND2_X1 U13050 ( .A1(n11121), .A2(n11120), .ZN(n15589) );
  XNOR2_X1 U13051 ( .A(n11122), .B(n7571), .ZN(n11132) );
  INV_X1 U13052 ( .A(n11132), .ZN(n16411) );
  INV_X1 U13053 ( .A(n16454), .ZN(n16387) );
  OAI22_X1 U13054 ( .A1(n7856), .A2(n16389), .B1(n11123), .B2(n15805), .ZN(
        n11127) );
  NAND2_X1 U13055 ( .A1(n11122), .A2(n13310), .ZN(n11124) );
  AOI21_X1 U13056 ( .B1(n11125), .B2(n11124), .A(n16558), .ZN(n11126) );
  AOI211_X1 U13057 ( .C1(n16411), .C2(n16387), .A(n11127), .B(n11126), .ZN(
        n16408) );
  OAI22_X1 U13058 ( .A1(n15812), .A2(n11130), .B1(n11129), .B2(n16395), .ZN(
        n11134) );
  NAND2_X1 U13059 ( .A1(n15812), .A2(n15519), .ZN(n15780) );
  INV_X1 U13060 ( .A(n11142), .ZN(n11131) );
  OAI211_X1 U13061 ( .C1(n7601), .C2(n13308), .A(n11131), .B(n15910), .ZN(
        n16407) );
  OR2_X1 U13062 ( .A1(n13028), .A2(n15519), .ZN(n12996) );
  INV_X1 U13063 ( .A(n12996), .ZN(n16399) );
  NAND2_X1 U13064 ( .A1(n15812), .A2(n16399), .ZN(n16547) );
  OAI22_X1 U13065 ( .A1(n15780), .A2(n16407), .B1(n16547), .B2(n11132), .ZN(
        n11133) );
  AOI211_X1 U13066 ( .C1(n16525), .C2(n13025), .A(n11134), .B(n11133), .ZN(
        n11135) );
  OAI21_X1 U13067 ( .B1(n16605), .B2(n16408), .A(n11135), .ZN(P1_U3292) );
  XNOR2_X1 U13068 ( .A(n11137), .B(n13313), .ZN(n16436) );
  OAI21_X1 U13069 ( .B1(n11139), .B2(n13313), .A(n11138), .ZN(n16439) );
  INV_X1 U13070 ( .A(n16395), .ZN(n16592) );
  AOI22_X1 U13071 ( .A1(n15812), .A2(n16431), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n16592), .ZN(n11140) );
  OAI21_X1 U13072 ( .B1(n11141), .B2(n15812), .A(n11140), .ZN(n11144) );
  OAI211_X1 U13073 ( .C1(n16434), .C2(n11142), .A(n15910), .B(n11174), .ZN(
        n16432) );
  OAI22_X1 U13074 ( .A1(n16434), .A2(n16595), .B1(n15780), .B2(n16432), .ZN(
        n11143) );
  AOI211_X1 U13075 ( .C1(n15711), .C2(n16439), .A(n11144), .B(n11143), .ZN(
        n11145) );
  OAI21_X1 U13076 ( .B1(n16597), .B2(n16436), .A(n11145), .ZN(P1_U3291) );
  AOI22_X1 U13077 ( .A1(n16036), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n11151) );
  NAND3_X1 U13078 ( .A1(n16382), .A2(n16374), .A3(n16376), .ZN(n11149) );
  OAI21_X1 U13079 ( .B1(P3_IR_REG_0__SCAN_IN), .B2(n11147), .A(n11146), .ZN(
        n11148) );
  NAND2_X1 U13080 ( .A1(n11149), .A2(n11148), .ZN(n11150) );
  OAI211_X1 U13081 ( .C1(n16367), .C2(n11152), .A(n11151), .B(n11150), .ZN(
        P3_U3182) );
  INV_X1 U13082 ( .A(n11153), .ZN(n11155) );
  NAND2_X1 U13083 ( .A1(n11155), .A2(n11154), .ZN(n11156) );
  XNOR2_X1 U13084 ( .A(n11157), .B(n11156), .ZN(n11161) );
  NAND2_X1 U13085 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n14798) );
  OAI21_X1 U13086 ( .B1(n14683), .B2(n12038), .A(n14798), .ZN(n11159) );
  OAI22_X1 U13087 ( .A1(n11465), .A2(n12029), .B1(n7947), .B2(n14705), .ZN(
        n11158) );
  AOI211_X1 U13088 ( .C1(n14702), .C2(n14727), .A(n11159), .B(n11158), .ZN(
        n11160) );
  OAI21_X1 U13089 ( .B1(n14686), .B2(n11161), .A(n11160), .ZN(P2_U3193) );
  OAI222_X1 U13090 ( .A1(n14150), .A2(n14424), .B1(P3_U3151), .B2(n13694), 
        .C1(n14154), .C2(n11162), .ZN(P3_U3276) );
  INV_X1 U13091 ( .A(n13127), .ZN(n11245) );
  AOI22_X1 U13092 ( .A1(n16102), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n11163), .ZN(n11164) );
  OAI21_X1 U13093 ( .B1(n11245), .B2(n15123), .A(n11164), .ZN(P2_U3310) );
  NAND2_X1 U13094 ( .A1(n11165), .A2(n16580), .ZN(n11166) );
  OR2_X1 U13095 ( .A1(n12926), .A2(n11166), .ZN(n11168) );
  NAND2_X1 U13096 ( .A1(n10734), .A2(n13967), .ZN(n11167) );
  AND2_X1 U13097 ( .A1(n11168), .A2(n11167), .ZN(n11246) );
  INV_X1 U13098 ( .A(n11246), .ZN(n11523) );
  INV_X1 U13099 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11169) );
  OAI22_X1 U13100 ( .A1(n14139), .A2(n11528), .B1(n16590), .B2(n11169), .ZN(
        n11170) );
  AOI21_X1 U13101 ( .B1(n11523), .B2(n16590), .A(n11170), .ZN(n11171) );
  INV_X1 U13102 ( .A(n11171), .ZN(P3_U3390) );
  XNOR2_X1 U13103 ( .A(n11172), .B(n13312), .ZN(n16453) );
  NAND2_X1 U13104 ( .A1(n11174), .A2(n11173), .ZN(n11175) );
  NAND3_X1 U13105 ( .A1(n11363), .A2(n15910), .A3(n11175), .ZN(n16451) );
  INV_X1 U13106 ( .A(n16451), .ZN(n11179) );
  MUX2_X1 U13107 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n11176), .S(n15812), .Z(
        n11178) );
  OAI22_X1 U13108 ( .A1(n16595), .A2(n16452), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n16395), .ZN(n11177) );
  AOI211_X1 U13109 ( .C1(n11179), .C2(n16601), .A(n11178), .B(n11177), .ZN(
        n11182) );
  XNOR2_X1 U13110 ( .A(n11180), .B(n13312), .ZN(n16457) );
  NAND2_X1 U13111 ( .A1(n16457), .A2(n15711), .ZN(n11181) );
  OAI211_X1 U13112 ( .C1(n16597), .C2(n16453), .A(n11182), .B(n11181), .ZN(
        P1_U3290) );
  MUX2_X1 U13113 ( .A(n11183), .B(P1_REG2_REG_5__SCAN_IN), .S(n16605), .Z(
        n11184) );
  INV_X1 U13114 ( .A(n11184), .ZN(n11189) );
  OAI22_X1 U13115 ( .A1(n16595), .A2(n13054), .B1(n16395), .B2(n11185), .ZN(
        n11186) );
  AOI21_X1 U13116 ( .B1(n11187), .B2(n16601), .A(n11186), .ZN(n11188) );
  OAI211_X1 U13117 ( .C1(n11190), .C2(n16547), .A(n11189), .B(n11188), .ZN(
        P1_U3288) );
  INV_X1 U13118 ( .A(n11191), .ZN(n11192) );
  XNOR2_X1 U13119 ( .A(n11500), .B(n11194), .ZN(n11195) );
  AOI21_X1 U13120 ( .B1(n11196), .B2(n11195), .A(n13480), .ZN(n11201) );
  AOI22_X1 U13121 ( .A1(n13589), .A2(n10734), .B1(n13607), .B2(n13566), .ZN(
        n11197) );
  OAI21_X1 U13122 ( .B1(n12798), .B2(n13582), .A(n11197), .ZN(n11198) );
  AOI21_X1 U13123 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n11199), .A(n11198), .ZN(
        n11200) );
  OAI21_X1 U13124 ( .B1(n11201), .B2(n13599), .A(n11200), .ZN(P3_U3177) );
  OAI21_X1 U13125 ( .B1(n11203), .B2(n13315), .A(n11202), .ZN(n11209) );
  INV_X1 U13126 ( .A(n11209), .ZN(n16494) );
  OAI22_X1 U13127 ( .A1(n11204), .A2(n15805), .B1(n11566), .B2(n16389), .ZN(
        n11208) );
  XNOR2_X1 U13128 ( .A(n11205), .B(n13059), .ZN(n11206) );
  NOR2_X1 U13129 ( .A1(n11206), .A2(n16558), .ZN(n11207) );
  AOI211_X1 U13130 ( .C1(n16387), .C2(n11209), .A(n11208), .B(n11207), .ZN(
        n16492) );
  MUX2_X1 U13131 ( .A(n11210), .B(n16492), .S(n15812), .Z(n11219) );
  INV_X1 U13132 ( .A(n11211), .ZN(n11214) );
  INV_X1 U13133 ( .A(n11212), .ZN(n11213) );
  AOI211_X1 U13134 ( .C1(n16489), .C2(n11214), .A(n15915), .B(n11213), .ZN(
        n16488) );
  OAI22_X1 U13135 ( .A1(n16595), .A2(n11216), .B1(n11215), .B2(n16395), .ZN(
        n11217) );
  AOI21_X1 U13136 ( .B1(n16488), .B2(n16601), .A(n11217), .ZN(n11218) );
  OAI211_X1 U13137 ( .C1(n16494), .C2(n16547), .A(n11219), .B(n11218), .ZN(
        P1_U3287) );
  INV_X1 U13138 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n12280) );
  MUX2_X1 U13139 ( .A(n12285), .B(n12280), .S(n7429), .Z(n11220) );
  NAND2_X1 U13140 ( .A1(n11220), .A2(n7908), .ZN(n11389) );
  OAI21_X1 U13141 ( .B1(n11220), .B2(n7908), .A(n11389), .ZN(n11225) );
  AOI21_X1 U13142 ( .B1(n11225), .B2(n11224), .A(n11397), .ZN(n11241) );
  XNOR2_X1 U13143 ( .A(n11386), .B(P3_REG2_REG_7__SCAN_IN), .ZN(n11239) );
  INV_X1 U13144 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11229) );
  OR2_X1 U13145 ( .A1(n11230), .A2(n11229), .ZN(n11231) );
  NAND2_X1 U13146 ( .A1(n11233), .A2(n12280), .ZN(n11234) );
  AOI21_X1 U13147 ( .B1(n11405), .B2(n11234), .A(n16374), .ZN(n11238) );
  INV_X1 U13148 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n11235) );
  NOR2_X1 U13149 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11235), .ZN(n13444) );
  AOI21_X1 U13150 ( .B1(n16036), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n13444), .ZN(
        n11236) );
  OAI21_X1 U13151 ( .B1(n16367), .B2(n11385), .A(n11236), .ZN(n11237) );
  AOI211_X1 U13152 ( .C1(n13712), .C2(n11239), .A(n11238), .B(n11237), .ZN(
        n11240) );
  OAI21_X1 U13153 ( .B1(n11241), .B2(n16376), .A(n11240), .ZN(P3_U3189) );
  NAND2_X1 U13154 ( .A1(n11242), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11243) );
  XNOR2_X1 U13155 ( .A(n11243), .B(n14606), .ZN(n13128) );
  OAI222_X1 U13156 ( .A1(n13128), .A2(P1_U3086), .B1(n15990), .B2(n11245), 
        .C1(n11244), .C2(n15992), .ZN(P1_U3338) );
  MUX2_X1 U13157 ( .A(n11246), .B(n9586), .S(n16585), .Z(n11247) );
  OAI21_X1 U13158 ( .B1(n11528), .B2(n14051), .A(n11247), .ZN(P3_U3459) );
  XNOR2_X1 U13159 ( .A(n11249), .B(n11248), .ZN(n11250) );
  INV_X1 U13160 ( .A(n16376), .ZN(n11900) );
  NAND2_X1 U13161 ( .A1(n11250), .A2(n11900), .ZN(n11265) );
  OAI21_X1 U13162 ( .B1(n11253), .B2(n11252), .A(n11251), .ZN(n11263) );
  INV_X1 U13163 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n16196) );
  NOR2_X1 U13164 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11254), .ZN(n11508) );
  INV_X1 U13165 ( .A(n11508), .ZN(n11255) );
  OAI21_X1 U13166 ( .B1(n16364), .B2(n16196), .A(n11255), .ZN(n11262) );
  INV_X1 U13167 ( .A(n11256), .ZN(n11258) );
  NAND3_X1 U13168 ( .A1(n11272), .A2(n11258), .A3(n11257), .ZN(n11259) );
  AOI21_X1 U13169 ( .B1(n11260), .B2(n11259), .A(n16374), .ZN(n11261) );
  AOI211_X1 U13170 ( .C1(n13712), .C2(n11263), .A(n11262), .B(n11261), .ZN(
        n11264) );
  OAI211_X1 U13171 ( .C1(n16367), .C2(n11266), .A(n11265), .B(n11264), .ZN(
        P3_U3186) );
  XOR2_X1 U13172 ( .A(n11267), .B(n11268), .Z(n11279) );
  XOR2_X1 U13173 ( .A(n11269), .B(P3_REG2_REG_3__SCAN_IN), .Z(n11275) );
  NOR2_X1 U13174 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14472), .ZN(n13482) );
  NAND2_X1 U13175 ( .A1(n11270), .A2(n16448), .ZN(n11271) );
  AOI21_X1 U13176 ( .B1(n11272), .B2(n11271), .A(n16374), .ZN(n11273) );
  AOI211_X1 U13177 ( .C1(n16036), .C2(P3_ADDR_REG_3__SCAN_IN), .A(n13482), .B(
        n11273), .ZN(n11274) );
  OAI21_X1 U13178 ( .B1(n11275), .B2(n16382), .A(n11274), .ZN(n11276) );
  AOI21_X1 U13179 ( .B1(n11277), .B2(n13707), .A(n11276), .ZN(n11278) );
  OAI21_X1 U13180 ( .B1(n11279), .B2(n16376), .A(n11278), .ZN(P3_U3185) );
  INV_X1 U13181 ( .A(n11280), .ZN(n11283) );
  INV_X1 U13182 ( .A(SI_20_), .ZN(n11282) );
  OAI222_X1 U13183 ( .A1(n14154), .A2(n11283), .B1(n14150), .B2(n11282), .C1(
        P3_U3151), .C2(n11281), .ZN(P3_U3275) );
  INV_X1 U13184 ( .A(n11286), .ZN(n11288) );
  OR2_X1 U13185 ( .A1(n11288), .A2(n11287), .ZN(n11289) );
  OR2_X1 U13186 ( .A1(n11290), .A2(n12973), .ZN(n11292) );
  AOI22_X1 U13187 ( .A1(n13155), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n13154), 
        .B2(n15462), .ZN(n11291) );
  NAND2_X1 U13188 ( .A1(n16526), .A2(n15255), .ZN(n11294) );
  NAND2_X1 U13189 ( .A1(n15377), .A2(n7432), .ZN(n11293) );
  NAND2_X1 U13190 ( .A1(n11294), .A2(n11293), .ZN(n11295) );
  XNOR2_X1 U13191 ( .A(n11295), .B(n15221), .ZN(n11298) );
  INV_X1 U13192 ( .A(n15377), .ZN(n11590) );
  NOR2_X1 U13193 ( .A1(n11590), .A2(n15223), .ZN(n11296) );
  AOI21_X1 U13194 ( .B1(n16526), .B2(n7432), .A(n11296), .ZN(n11297) );
  NAND2_X1 U13195 ( .A1(n11298), .A2(n11297), .ZN(n11414) );
  OR2_X1 U13196 ( .A1(n11298), .A2(n11297), .ZN(n11299) );
  NAND2_X1 U13197 ( .A1(n11414), .A2(n11299), .ZN(n11301) );
  INV_X1 U13198 ( .A(n11415), .ZN(n11300) );
  AOI21_X1 U13199 ( .B1(n11302), .B2(n11301), .A(n11300), .ZN(n11314) );
  NAND2_X1 U13200 ( .A1(n13170), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n11310) );
  OR2_X1 U13201 ( .A1(n13256), .A2(n11303), .ZN(n11309) );
  AND2_X1 U13202 ( .A1(n11305), .A2(n11304), .ZN(n11306) );
  OR2_X1 U13203 ( .A1(n11306), .A2(n11429), .ZN(n16543) );
  OR2_X1 U13204 ( .A1(n13282), .A2(n16543), .ZN(n11308) );
  OR2_X1 U13205 ( .A1(n13284), .A2(n11823), .ZN(n11307) );
  NAND4_X1 U13206 ( .A1(n11310), .A2(n11309), .A3(n11308), .A4(n11307), .ZN(
        n15376) );
  INV_X1 U13207 ( .A(n15376), .ZN(n11592) );
  OAI22_X1 U13208 ( .A1(n11566), .A2(n15805), .B1(n11592), .B2(n16389), .ZN(
        n11571) );
  NAND2_X1 U13209 ( .A1(n15277), .A2(n11571), .ZN(n11311) );
  NAND2_X1 U13210 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n15460) );
  OAI211_X1 U13211 ( .C1(n15360), .C2(n16523), .A(n11311), .B(n15460), .ZN(
        n11312) );
  AOI21_X1 U13212 ( .B1(n16526), .B2(n15365), .A(n11312), .ZN(n11313) );
  OAI21_X1 U13213 ( .B1(n11314), .B2(n15367), .A(n11313), .ZN(P1_U3221) );
  INV_X1 U13214 ( .A(n11315), .ZN(n11316) );
  AND3_X1 U13215 ( .A1(n16040), .A2(n11316), .A3(n16039), .ZN(n11317) );
  NAND2_X1 U13216 ( .A1(n11318), .A2(n11317), .ZN(n11787) );
  NAND2_X1 U13217 ( .A1(n11319), .A2(n11851), .ZN(n11320) );
  NOR2_X1 U13218 ( .A1(n14922), .A2(n10594), .ZN(n11321) );
  AOI211_X1 U13219 ( .C1(n11324), .C2(n11323), .A(n11322), .B(n11321), .ZN(
        n11325) );
  NOR2_X1 U13220 ( .A1(n11325), .A2(n14992), .ZN(n11326) );
  AOI21_X1 U13221 ( .B1(n16522), .B2(P2_REG2_REG_0__SCAN_IN), .A(n11326), .ZN(
        n11327) );
  OAI21_X1 U13222 ( .B1(n11328), .B2(n14829), .A(n11327), .ZN(P2_U3265) );
  NOR2_X1 U13223 ( .A1(n16595), .A2(n11329), .ZN(n11335) );
  MUX2_X1 U13224 ( .A(n11331), .B(n11330), .S(n15812), .Z(n11332) );
  OAI21_X1 U13225 ( .B1(n16395), .B2(n11333), .A(n11332), .ZN(n11334) );
  AOI211_X1 U13226 ( .C1(n11336), .C2(n16601), .A(n11335), .B(n11334), .ZN(
        n11339) );
  INV_X1 U13227 ( .A(n16597), .ZN(n15818) );
  NAND2_X1 U13228 ( .A1(n11337), .A2(n15818), .ZN(n11338) );
  OAI211_X1 U13229 ( .C1(n11340), .C2(n15821), .A(n11339), .B(n11338), .ZN(
        P1_U3286) );
  NAND2_X1 U13230 ( .A1(n11802), .A2(n14731), .ZN(n11342) );
  NAND2_X1 U13231 ( .A1(n11343), .A2(n11353), .ZN(n11545) );
  OAI21_X1 U13232 ( .B1(n11343), .B2(n11353), .A(n11545), .ZN(n16518) );
  INV_X1 U13233 ( .A(n16518), .ZN(n11358) );
  AND2_X1 U13234 ( .A1(n11344), .A2(n11802), .ZN(n11345) );
  NAND2_X1 U13235 ( .A1(n11347), .A2(n14731), .ZN(n11348) );
  INV_X1 U13236 ( .A(n11918), .ZN(n11923) );
  NAND2_X1 U13237 ( .A1(n11934), .A2(n11350), .ZN(n11352) );
  INV_X1 U13238 ( .A(n11353), .ZN(n11351) );
  NAND3_X1 U13239 ( .A1(n11920), .A2(n11353), .A3(n11352), .ZN(n11354) );
  NAND2_X1 U13240 ( .A1(n11549), .A2(n11354), .ZN(n11355) );
  AOI222_X1 U13241 ( .A1(n14981), .A2(n11355), .B1(n14728), .B2(n14913), .C1(
        n14730), .C2(n14911), .ZN(n16505) );
  INV_X1 U13242 ( .A(n11928), .ZN(n11356) );
  AOI211_X1 U13243 ( .C1(n11548), .C2(n11356), .A(n14986), .B(n7948), .ZN(
        n16509) );
  AOI21_X1 U13244 ( .B1(n15079), .B2(n11548), .A(n16509), .ZN(n11357) );
  OAI211_X1 U13245 ( .C1(n15082), .C2(n11358), .A(n16505), .B(n11357), .ZN(
        n11373) );
  NAND2_X1 U13246 ( .A1(n11373), .A2(n7433), .ZN(n11359) );
  OAI21_X1 U13247 ( .B1(n7433), .B2(n10295), .A(n11359), .ZN(P2_U3506) );
  XNOR2_X1 U13248 ( .A(n11362), .B(n15381), .ZN(n13317) );
  XNOR2_X1 U13249 ( .A(n11360), .B(n13317), .ZN(n11361) );
  AOI222_X1 U13250 ( .A1(n16458), .A2(n11361), .B1(n15380), .B2(n15789), .C1(
        n15382), .C2(n15787), .ZN(n16464) );
  NAND2_X1 U13251 ( .A1(n11363), .A2(n11362), .ZN(n11364) );
  NAND2_X1 U13252 ( .A1(n11364), .A2(n15910), .ZN(n11365) );
  NOR2_X1 U13253 ( .A1(n11366), .A2(n11365), .ZN(n16461) );
  OAI22_X1 U13254 ( .A1(n15812), .A2(n10528), .B1(n11367), .B2(n16395), .ZN(
        n11369) );
  NOR2_X1 U13255 ( .A1(n16595), .A2(n16463), .ZN(n11368) );
  AOI211_X1 U13256 ( .C1(n16461), .C2(n16601), .A(n11369), .B(n11368), .ZN(
        n11372) );
  XOR2_X1 U13257 ( .A(n13317), .B(n11370), .Z(n16467) );
  NAND2_X1 U13258 ( .A1(n16467), .A2(n15818), .ZN(n11371) );
  OAI211_X1 U13259 ( .C1(n16464), .C2(n16605), .A(n11372), .B(n11371), .ZN(
        P1_U3289) );
  NAND2_X1 U13260 ( .A1(n11373), .A2(n15102), .ZN(n11374) );
  OAI21_X1 U13261 ( .B1(n15102), .B2(n8699), .A(n11374), .ZN(P2_U3451) );
  INV_X1 U13262 ( .A(n11375), .ZN(n11376) );
  AOI21_X1 U13263 ( .B1(n11378), .B2(n11377), .A(n11376), .ZN(n11382) );
  AOI22_X1 U13264 ( .A1(n14701), .A2(n14728), .B1(n14702), .B2(n14726), .ZN(
        n11379) );
  NAND2_X1 U13265 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n16154) );
  OAI211_X1 U13266 ( .C1(n12097), .C2(n14683), .A(n11379), .B(n16154), .ZN(
        n11380) );
  AOI21_X1 U13267 ( .B1(n12095), .B2(n14691), .A(n11380), .ZN(n11381) );
  OAI21_X1 U13268 ( .B1(n11382), .B2(n14686), .A(n11381), .ZN(P2_U3203) );
  MUX2_X1 U13269 ( .A(P3_REG2_REG_8__SCAN_IN), .B(n11390), .S(n11665), .Z(
        n11388) );
  INV_X1 U13270 ( .A(n11383), .ZN(n11384) );
  NOR2_X1 U13271 ( .A1(n11387), .A2(n11388), .ZN(n11662) );
  AOI21_X1 U13272 ( .B1(n11388), .B2(n11387), .A(n11662), .ZN(n11411) );
  INV_X1 U13273 ( .A(n11389), .ZN(n11396) );
  INV_X1 U13274 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n12249) );
  MUX2_X1 U13275 ( .A(n11390), .B(n12249), .S(n7429), .Z(n11391) );
  NAND2_X1 U13276 ( .A1(n11391), .A2(n11665), .ZN(n11680) );
  INV_X1 U13277 ( .A(n11391), .ZN(n11393) );
  NAND2_X1 U13278 ( .A1(n11393), .A2(n11392), .ZN(n11394) );
  AND2_X1 U13279 ( .A1(n11680), .A2(n11394), .ZN(n11395) );
  INV_X1 U13280 ( .A(n11681), .ZN(n11399) );
  NOR3_X1 U13281 ( .A1(n11397), .A2(n11396), .A3(n11395), .ZN(n11398) );
  OAI21_X1 U13282 ( .B1(n11399), .B2(n11398), .A(n11900), .ZN(n11410) );
  INV_X1 U13283 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n16246) );
  NOR2_X1 U13284 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14273), .ZN(n12393) );
  INV_X1 U13285 ( .A(n12393), .ZN(n11400) );
  OAI21_X1 U13286 ( .B1(n16364), .B2(n16246), .A(n11400), .ZN(n11408) );
  NAND2_X1 U13287 ( .A1(n11405), .A2(n11403), .ZN(n11401) );
  MUX2_X1 U13288 ( .A(n12249), .B(P3_REG1_REG_8__SCAN_IN), .S(n11665), .Z(
        n11402) );
  NAND2_X1 U13289 ( .A1(n11401), .A2(n11402), .ZN(n11667) );
  INV_X1 U13290 ( .A(n11402), .ZN(n11404) );
  NAND3_X1 U13291 ( .A1(n11405), .A2(n11404), .A3(n11403), .ZN(n11406) );
  AOI21_X1 U13292 ( .B1(n11667), .B2(n11406), .A(n16374), .ZN(n11407) );
  AOI211_X1 U13293 ( .C1(n13707), .C2(n11665), .A(n11408), .B(n11407), .ZN(
        n11409) );
  OAI211_X1 U13294 ( .C1(n11411), .C2(n16382), .A(n11410), .B(n11409), .ZN(
        P3_U3190) );
  INV_X1 U13295 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n11413) );
  NAND2_X1 U13296 ( .A1(n13421), .A2(n11644), .ZN(n11412) );
  OAI21_X1 U13297 ( .B1(P3_U3897), .B2(n11413), .A(n11412), .ZN(P3_U3517) );
  NAND2_X1 U13298 ( .A1(n11416), .A2(n13289), .ZN(n11418) );
  AOI22_X1 U13299 ( .A1(n13155), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n15478), 
        .B2(n13154), .ZN(n11417) );
  NAND2_X1 U13300 ( .A1(n13078), .A2(n15255), .ZN(n11420) );
  NAND2_X1 U13301 ( .A1(n15376), .A2(n7432), .ZN(n11419) );
  NAND2_X1 U13302 ( .A1(n11420), .A2(n11419), .ZN(n11421) );
  XNOR2_X1 U13303 ( .A(n11421), .B(n15253), .ZN(n11424) );
  NAND2_X1 U13304 ( .A1(n13078), .A2(n7432), .ZN(n11423) );
  OR2_X1 U13305 ( .A1(n11592), .A2(n15223), .ZN(n11422) );
  NAND2_X1 U13306 ( .A1(n11423), .A2(n11422), .ZN(n11425) );
  NAND2_X1 U13307 ( .A1(n11424), .A2(n11425), .ZN(n11611) );
  INV_X1 U13308 ( .A(n11424), .ZN(n11427) );
  INV_X1 U13309 ( .A(n11425), .ZN(n11426) );
  NAND2_X1 U13310 ( .A1(n11427), .A2(n11426), .ZN(n11613) );
  NAND2_X1 U13311 ( .A1(n11611), .A2(n11613), .ZN(n11428) );
  XNOR2_X1 U13312 ( .A(n11612), .B(n11428), .ZN(n11440) );
  NAND2_X1 U13313 ( .A1(n13170), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n11434) );
  OR2_X1 U13314 ( .A1(n13256), .A2(n11595), .ZN(n11433) );
  NOR2_X1 U13315 ( .A1(n11429), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11430) );
  OR2_X1 U13316 ( .A1(n11598), .A2(n11430), .ZN(n11622) );
  OR2_X1 U13317 ( .A1(n13282), .A2(n11622), .ZN(n11432) );
  OR2_X1 U13318 ( .A1(n13284), .A2(n16566), .ZN(n11431) );
  NAND4_X1 U13319 ( .A1(n11434), .A2(n11433), .A3(n11432), .A4(n11431), .ZN(
        n15375) );
  NAND2_X1 U13320 ( .A1(n15789), .A2(n15375), .ZN(n11436) );
  NAND2_X1 U13321 ( .A1(n15787), .A2(n15377), .ZN(n11435) );
  NAND2_X1 U13322 ( .A1(n11436), .A2(n11435), .ZN(n11813) );
  NAND2_X1 U13323 ( .A1(n15277), .A2(n11813), .ZN(n11437) );
  NAND2_X1 U13324 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n15475) );
  OAI211_X1 U13325 ( .C1(n15360), .C2(n16543), .A(n11437), .B(n15475), .ZN(
        n11438) );
  AOI21_X1 U13326 ( .B1(n13078), .B2(n15365), .A(n11438), .ZN(n11439) );
  OAI21_X1 U13327 ( .B1(n11440), .B2(n15367), .A(n11439), .ZN(P1_U3231) );
  INV_X1 U13328 ( .A(n11441), .ZN(n11444) );
  INV_X1 U13329 ( .A(SI_21_), .ZN(n11443) );
  OAI222_X1 U13330 ( .A1(n14154), .A2(n11444), .B1(n14150), .B2(n11443), .C1(
        P3_U3151), .C2(n11442), .ZN(P3_U3274) );
  INV_X1 U13331 ( .A(n11445), .ZN(n12000) );
  NAND2_X1 U13332 ( .A1(n12000), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11448) );
  INV_X1 U13333 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11446) );
  MUX2_X1 U13334 ( .A(n11446), .B(P1_REG2_REG_14__SCAN_IN), .S(n12313), .Z(
        n11447) );
  AOI21_X1 U13335 ( .B1(n11449), .B2(n11448), .A(n11447), .ZN(n11486) );
  INV_X1 U13336 ( .A(n11486), .ZN(n11451) );
  NAND3_X1 U13337 ( .A1(n11449), .A2(n11448), .A3(n11447), .ZN(n11450) );
  NAND3_X1 U13338 ( .A1(n11451), .A2(n15516), .A3(n11450), .ZN(n11457) );
  NAND2_X1 U13339 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n12522)
         );
  XOR2_X1 U13340 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n11485), .Z(n11453) );
  NAND2_X1 U13341 ( .A1(n15517), .A2(n11453), .ZN(n11454) );
  NAND2_X1 U13342 ( .A1(n12522), .A2(n11454), .ZN(n11455) );
  AOI21_X1 U13343 ( .B1(n16162), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n11455), 
        .ZN(n11456) );
  OAI211_X1 U13344 ( .C1(n15511), .C2(n11458), .A(n11457), .B(n11456), .ZN(
        P1_U3257) );
  INV_X1 U13345 ( .A(n12151), .ZN(n16573) );
  OAI21_X1 U13346 ( .B1(n11461), .B2(n11460), .A(n11459), .ZN(n11462) );
  NAND2_X1 U13347 ( .A1(n11462), .A2(n14707), .ZN(n11470) );
  INV_X1 U13348 ( .A(n12148), .ZN(n11468) );
  OAI22_X1 U13349 ( .A1(n12065), .A2(n11465), .B1(n11464), .B2(n11463), .ZN(
        n11466) );
  AOI211_X1 U13350 ( .C1(n11468), .C2(n14700), .A(n11467), .B(n11466), .ZN(
        n11469) );
  OAI211_X1 U13351 ( .C1(n16573), .C2(n14705), .A(n11470), .B(n11469), .ZN(
        P2_U3189) );
  INV_X1 U13352 ( .A(n13135), .ZN(n11494) );
  NAND2_X1 U13353 ( .A1(n11471), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11472) );
  XNOR2_X1 U13354 ( .A(n11472), .B(P1_IR_REG_18__SCAN_IN), .ZN(n15507) );
  INV_X1 U13355 ( .A(n15507), .ZN(n12585) );
  OAI222_X1 U13356 ( .A1(n15987), .A2(n11473), .B1(n15990), .B2(n11494), .C1(
        P1_U3086), .C2(n12585), .ZN(P1_U3337) );
  XNOR2_X1 U13357 ( .A(n11474), .B(n7578), .ZN(n11690) );
  NAND2_X1 U13358 ( .A1(n11942), .A2(n11475), .ZN(n11476) );
  XNOR2_X1 U13359 ( .A(n9995), .B(n11476), .ZN(n11478) );
  AOI22_X1 U13360 ( .A1(n13954), .A2(n13607), .B1(n12163), .B2(n13967), .ZN(
        n11477) );
  OAI21_X1 U13361 ( .B1(n11478), .B2(n13878), .A(n11477), .ZN(n11479) );
  AOI21_X1 U13362 ( .B1(n11690), .B2(n14052), .A(n11479), .ZN(n11688) );
  NAND2_X1 U13363 ( .A1(n16590), .A2(n16485), .ZN(n14109) );
  OAI22_X1 U13364 ( .A1(n14139), .A2(n8016), .B1(n16590), .B2(n11480), .ZN(
        n11481) );
  AOI21_X1 U13365 ( .B1(n11690), .B2(n14134), .A(n11481), .ZN(n11482) );
  OAI21_X1 U13366 ( .B1(n11688), .B2(n16588), .A(n11482), .ZN(P3_U3402) );
  INV_X1 U13367 ( .A(n11483), .ZN(n11484) );
  AOI22_X1 U13368 ( .A1(n11485), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n12313), 
        .B2(n11484), .ZN(n12214) );
  XNOR2_X1 U13369 ( .A(n12212), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n11493) );
  INV_X1 U13370 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n16315) );
  NAND2_X1 U13371 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15357)
         );
  OAI21_X1 U13372 ( .B1(n15524), .B2(n16315), .A(n15357), .ZN(n11491) );
  AOI21_X1 U13373 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n12313), .A(n11486), 
        .ZN(n11487) );
  NAND2_X1 U13374 ( .A1(n11487), .A2(n12213), .ZN(n12209) );
  OAI21_X1 U13375 ( .B1(n11487), .B2(n12213), .A(n12209), .ZN(n11488) );
  NOR2_X1 U13376 ( .A1(n11488), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n12208) );
  AOI21_X1 U13377 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n11488), .A(n12208), 
        .ZN(n11489) );
  NOR2_X1 U13378 ( .A1(n11489), .A2(n15512), .ZN(n11490) );
  AOI211_X1 U13379 ( .C1(n15477), .C2(n12403), .A(n11491), .B(n11490), .ZN(
        n11492) );
  OAI21_X1 U13380 ( .B1(n11493), .B2(n15398), .A(n11492), .ZN(P1_U3258) );
  INV_X1 U13381 ( .A(n16115), .ZN(n11847) );
  OAI222_X1 U13382 ( .A1(n15133), .A2(n11495), .B1(n11847), .B2(P2_U3088), 
        .C1(n15123), .C2(n11494), .ZN(P2_U3309) );
  INV_X1 U13383 ( .A(n11496), .ZN(n11498) );
  OAI22_X1 U13384 ( .A1(n12963), .A2(P3_U3151), .B1(SI_22_), .B2(n14150), .ZN(
        n11497) );
  AOI21_X1 U13385 ( .B1(n11498), .B2(n11702), .A(n11497), .ZN(P3_U3273) );
  INV_X1 U13386 ( .A(n11640), .ZN(n11511) );
  XNOR2_X1 U13387 ( .A(n13484), .B(n11499), .ZN(n11502) );
  INV_X1 U13388 ( .A(n11502), .ZN(n11503) );
  NOR2_X1 U13389 ( .A1(n11500), .A2(n13483), .ZN(n13479) );
  XNOR2_X1 U13390 ( .A(n11502), .B(n11501), .ZN(n13478) );
  XNOR2_X1 U13391 ( .A(n11689), .B(n13425), .ZN(n11504) );
  NOR2_X1 U13392 ( .A1(n11504), .A2(n13485), .ZN(n11707) );
  AOI21_X1 U13393 ( .B1(n13485), .B2(n11504), .A(n11707), .ZN(n11505) );
  OAI21_X1 U13394 ( .B1(n7565), .B2(n11505), .A(n11709), .ZN(n11506) );
  NAND2_X1 U13395 ( .A1(n11506), .A2(n13576), .ZN(n11510) );
  OAI22_X1 U13396 ( .A1(n13582), .A2(n8016), .B1(n11754), .B2(n13593), .ZN(
        n11507) );
  AOI211_X1 U13397 ( .C1(n13589), .C2(n13607), .A(n11508), .B(n11507), .ZN(
        n11509) );
  OAI211_X1 U13398 ( .C1(n11511), .C2(n13448), .A(n11510), .B(n11509), .ZN(
        P3_U3170) );
  NAND2_X1 U13399 ( .A1(n13606), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n11512) );
  OAI21_X1 U13400 ( .B1(n12913), .B2(n13606), .A(n11512), .ZN(P3_U3521) );
  OR2_X1 U13401 ( .A1(n11516), .A2(n14141), .ZN(n11519) );
  NAND2_X1 U13402 ( .A1(n11514), .A2(n11513), .ZN(n11515) );
  NAND2_X1 U13403 ( .A1(n11516), .A2(n11515), .ZN(n11518) );
  NAND3_X1 U13404 ( .A1(n11519), .A2(n11518), .A3(n11517), .ZN(n11524) );
  INV_X1 U13405 ( .A(n11524), .ZN(n11521) );
  NOR2_X1 U13406 ( .A1(n12920), .A2(n16580), .ZN(n11520) );
  AOI21_X1 U13407 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n13980), .A(n11523), .ZN(
        n11526) );
  MUX2_X1 U13408 ( .A(n11526), .B(n11525), .S(n13910), .Z(n11527) );
  OAI21_X1 U13409 ( .B1(n11528), .B2(n13940), .A(n11527), .ZN(P3_U3233) );
  NOR2_X1 U13410 ( .A1(n11529), .A2(n16580), .ZN(n16403) );
  OAI21_X1 U13411 ( .B1(n12922), .B2(n11031), .A(n11530), .ZN(n11531) );
  NAND2_X1 U13412 ( .A1(n11531), .A2(n13973), .ZN(n11533) );
  AOI22_X1 U13413 ( .A1(n13967), .A2(n13483), .B1(n10636), .B2(n13954), .ZN(
        n11532) );
  NAND2_X1 U13414 ( .A1(n11533), .A2(n11532), .ZN(n16402) );
  AOI21_X1 U13415 ( .B1(n16403), .B2(n11534), .A(n16402), .ZN(n11535) );
  MUX2_X1 U13416 ( .A(n11536), .B(n11535), .S(n13977), .Z(n11540) );
  XNOR2_X1 U13417 ( .A(n11537), .B(n12922), .ZN(n16404) );
  AND2_X1 U13418 ( .A1(n12920), .A2(n12789), .ZN(n11635) );
  OR2_X1 U13419 ( .A1(n14052), .A2(n11635), .ZN(n11538) );
  AOI22_X1 U13420 ( .A1(n16404), .A2(n13942), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n13980), .ZN(n11539) );
  NAND2_X1 U13421 ( .A1(n11540), .A2(n11539), .ZN(P3_U3232) );
  INV_X1 U13422 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n11543) );
  INV_X1 U13423 ( .A(n13754), .ZN(n11541) );
  NAND2_X1 U13424 ( .A1(n11541), .A2(n11644), .ZN(n11542) );
  OAI21_X1 U13425 ( .B1(P3_U3897), .B2(n11543), .A(n11542), .ZN(P3_U3519) );
  OR2_X1 U13426 ( .A1(n11548), .A2(n14729), .ZN(n11544) );
  NAND2_X1 U13427 ( .A1(n12034), .A2(n14728), .ZN(n11546) );
  INV_X1 U13428 ( .A(n12069), .ZN(n11547) );
  XNOR2_X1 U13429 ( .A(n12070), .B(n11547), .ZN(n12102) );
  INV_X1 U13430 ( .A(n12102), .ZN(n11557) );
  NAND2_X1 U13431 ( .A1(n11548), .A2(n12029), .ZN(n12024) );
  NAND2_X1 U13432 ( .A1(n11550), .A2(n12033), .ZN(n12027) );
  NAND2_X1 U13433 ( .A1(n12034), .A2(n11551), .ZN(n11552) );
  NAND2_X1 U13434 ( .A1(n12027), .A2(n11552), .ZN(n12064) );
  XNOR2_X1 U13435 ( .A(n12064), .B(n12069), .ZN(n11554) );
  AOI22_X1 U13436 ( .A1(n14911), .A2(n14728), .B1(n14726), .B2(n14913), .ZN(
        n11553) );
  OAI21_X1 U13437 ( .B1(n11554), .B2(n14949), .A(n11553), .ZN(n11555) );
  AOI21_X1 U13438 ( .B1(n16507), .B2(n12102), .A(n11555), .ZN(n12105) );
  AOI211_X1 U13439 ( .C1(n12095), .C2(n12036), .A(n14986), .B(n12147), .ZN(
        n12101) );
  AOI21_X1 U13440 ( .B1(n15079), .B2(n12095), .A(n12101), .ZN(n11556) );
  OAI211_X1 U13441 ( .C1(n11557), .C2(n10450), .A(n12105), .B(n11556), .ZN(
        n11559) );
  NAND2_X1 U13442 ( .A1(n11559), .A2(n7433), .ZN(n11558) );
  OAI21_X1 U13443 ( .B1(n7433), .B2(n10302), .A(n11558), .ZN(P2_U3508) );
  NAND2_X1 U13444 ( .A1(n11559), .A2(n15102), .ZN(n11560) );
  OAI21_X1 U13445 ( .B1(n15102), .B2(n8738), .A(n11560), .ZN(P2_U3457) );
  INV_X1 U13446 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n11578) );
  OR2_X1 U13447 ( .A1(n13065), .A2(n15378), .ZN(n11561) );
  XNOR2_X1 U13448 ( .A(n16526), .B(n15377), .ZN(n13320) );
  NAND2_X1 U13449 ( .A1(n11564), .A2(n13320), .ZN(n11565) );
  AND2_X1 U13450 ( .A1(n11583), .A2(n11565), .ZN(n16529) );
  INV_X1 U13451 ( .A(n16529), .ZN(n11576) );
  NAND2_X1 U13452 ( .A1(n13065), .A2(n11566), .ZN(n11567) );
  AOI211_X1 U13453 ( .C1(n11563), .C2(n11569), .A(n16558), .B(n7566), .ZN(
        n11570) );
  AOI211_X1 U13454 ( .C1(n16387), .C2(n16529), .A(n11571), .B(n11570), .ZN(
        n16532) );
  NAND2_X1 U13455 ( .A1(n11572), .A2(n16526), .ZN(n11573) );
  NAND2_X1 U13456 ( .A1(n11573), .A2(n15910), .ZN(n11574) );
  NOR2_X1 U13457 ( .A1(n11815), .A2(n11574), .ZN(n16527) );
  AOI21_X1 U13458 ( .B1(n16490), .B2(n16526), .A(n16527), .ZN(n11575) );
  OAI211_X1 U13459 ( .C1(n16493), .C2(n11576), .A(n16532), .B(n11575), .ZN(
        n11579) );
  NAND2_X1 U13460 ( .A1(n11579), .A2(n16570), .ZN(n11577) );
  OAI21_X1 U13461 ( .B1(n16570), .B2(n11578), .A(n11577), .ZN(P1_U3483) );
  NAND2_X1 U13462 ( .A1(n11579), .A2(n16469), .ZN(n11580) );
  OAI21_X1 U13463 ( .B1(n16469), .B2(n11581), .A(n11580), .ZN(P1_U3536) );
  NAND2_X1 U13464 ( .A1(n16526), .A2(n15377), .ZN(n11582) );
  XNOR2_X1 U13465 ( .A(n13078), .B(n11592), .ZN(n13322) );
  OR2_X1 U13466 ( .A1(n13078), .A2(n15376), .ZN(n11584) );
  NAND2_X1 U13467 ( .A1(n11585), .A2(n13289), .ZN(n11587) );
  AOI22_X1 U13468 ( .A1(n15492), .A2(n13154), .B1(n13155), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n11586) );
  XNOR2_X1 U13469 ( .A(n13082), .B(n15375), .ZN(n13323) );
  INV_X1 U13470 ( .A(n13323), .ZN(n11588) );
  OAI21_X1 U13471 ( .B1(n11589), .B2(n11588), .A(n11861), .ZN(n16563) );
  INV_X1 U13472 ( .A(n16563), .ZN(n11610) );
  OR2_X1 U13473 ( .A1(n16526), .A2(n11590), .ZN(n11591) );
  NAND2_X1 U13474 ( .A1(n13078), .A2(n11592), .ZN(n11593) );
  INV_X1 U13475 ( .A(n11870), .ZN(n16559) );
  NOR2_X1 U13476 ( .A1(n11594), .A2(n13323), .ZN(n16560) );
  OR3_X1 U13477 ( .A1(n16559), .A2(n16560), .A3(n15821), .ZN(n11609) );
  NAND2_X1 U13478 ( .A1(n15787), .A2(n15376), .ZN(n16554) );
  MUX2_X1 U13479 ( .A(n11595), .B(n16554), .S(n15812), .Z(n11596) );
  OAI21_X1 U13480 ( .B1(n16395), .B2(n11622), .A(n11596), .ZN(n11607) );
  INV_X1 U13481 ( .A(n13078), .ZN(n16546) );
  INV_X1 U13482 ( .A(n11816), .ZN(n11597) );
  AOI21_X1 U13483 ( .B1(n11597), .B2(n13082), .A(n15915), .ZN(n11605) );
  INV_X1 U13484 ( .A(n13082), .ZN(n16557) );
  NAND2_X1 U13485 ( .A1(n13170), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n11604) );
  OR2_X1 U13486 ( .A1(n13256), .A2(n10556), .ZN(n11603) );
  OR2_X1 U13487 ( .A1(n11598), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n11599) );
  NAND2_X1 U13488 ( .A1(n11871), .A2(n11599), .ZN(n16591) );
  OR2_X1 U13489 ( .A1(n13282), .A2(n16591), .ZN(n11602) );
  OR2_X1 U13490 ( .A1(n13284), .A2(n11600), .ZN(n11601) );
  NAND4_X1 U13491 ( .A1(n11604), .A2(n11603), .A3(n11602), .A4(n11601), .ZN(
        n15374) );
  AOI22_X1 U13492 ( .A1(n11605), .A2(n7563), .B1(n15789), .B2(n15374), .ZN(
        n16555) );
  NOR2_X1 U13493 ( .A1(n16555), .A2(n15780), .ZN(n11606) );
  AOI211_X1 U13494 ( .C1(n16525), .C2(n13082), .A(n11607), .B(n11606), .ZN(
        n11608) );
  OAI211_X1 U13495 ( .C1(n11610), .C2(n16597), .A(n11609), .B(n11608), .ZN(
        P1_U3283) );
  NAND2_X1 U13496 ( .A1(n13082), .A2(n15255), .ZN(n11615) );
  NAND2_X1 U13497 ( .A1(n15375), .A2(n7432), .ZN(n11614) );
  NAND2_X1 U13498 ( .A1(n11615), .A2(n11614), .ZN(n11616) );
  XNOR2_X1 U13499 ( .A(n11616), .B(n15221), .ZN(n12053) );
  INV_X1 U13500 ( .A(n15375), .ZN(n11868) );
  NOR2_X1 U13501 ( .A1(n11868), .A2(n15223), .ZN(n11617) );
  AOI21_X1 U13502 ( .B1(n13082), .B2(n7432), .A(n11617), .ZN(n12052) );
  XNOR2_X1 U13503 ( .A(n12053), .B(n12052), .ZN(n11619) );
  AOI21_X1 U13504 ( .B1(n11618), .B2(n11619), .A(n15367), .ZN(n11621) );
  NAND2_X1 U13505 ( .A1(n11621), .A2(n12055), .ZN(n11625) );
  INV_X1 U13506 ( .A(n15359), .ZN(n15337) );
  AND2_X1 U13507 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n15491) );
  INV_X1 U13508 ( .A(n15374), .ZN(n12050) );
  OAI22_X1 U13509 ( .A1(n15362), .A2(n12050), .B1(n11622), .B2(n15360), .ZN(
        n11623) );
  AOI211_X1 U13510 ( .C1(n15337), .C2(n15376), .A(n15491), .B(n11623), .ZN(
        n11624) );
  OAI211_X1 U13511 ( .C1(n16557), .C2(n15340), .A(n11625), .B(n11624), .ZN(
        P1_U3217) );
  INV_X1 U13512 ( .A(n12792), .ZN(n11628) );
  INV_X1 U13513 ( .A(n11626), .ZN(n11627) );
  AOI21_X1 U13514 ( .B1(n11628), .B2(n11630), .A(n11627), .ZN(n11634) );
  AOI22_X1 U13515 ( .A1(n13485), .A2(n13967), .B1(n13954), .B2(n13483), .ZN(
        n11633) );
  AND2_X1 U13516 ( .A1(n11652), .A2(n11629), .ZN(n11631) );
  OAI211_X1 U13517 ( .C1(n11631), .C2(n11630), .A(n11942), .B(n13973), .ZN(
        n11632) );
  OAI211_X1 U13518 ( .C1(n11634), .C2(n14015), .A(n11633), .B(n11632), .ZN(
        n16445) );
  INV_X1 U13519 ( .A(n16445), .ZN(n11639) );
  INV_X1 U13520 ( .A(n11634), .ZN(n16447) );
  INV_X2 U13521 ( .A(n13958), .ZN(n13977) );
  INV_X1 U13522 ( .A(n13984), .ZN(n13846) );
  AOI22_X1 U13523 ( .A1(n13981), .A2(n13484), .B1(n13980), .B2(n14472), .ZN(
        n11636) );
  OAI21_X1 U13524 ( .B1(n9621), .B2(n13977), .A(n11636), .ZN(n11637) );
  AOI21_X1 U13525 ( .B1(n16447), .B2(n13846), .A(n11637), .ZN(n11638) );
  OAI21_X1 U13526 ( .B1(n11639), .B2(n13958), .A(n11638), .ZN(P3_U3230) );
  AOI22_X1 U13527 ( .A1(n13981), .A2(n11689), .B1(n13980), .B2(n11640), .ZN(
        n11641) );
  OAI21_X1 U13528 ( .B1(n10941), .B2(n13977), .A(n11641), .ZN(n11642) );
  AOI21_X1 U13529 ( .B1(n11690), .B2(n13846), .A(n11642), .ZN(n11643) );
  OAI21_X1 U13530 ( .B1(n11688), .B2(n13958), .A(n11643), .ZN(P3_U3229) );
  INV_X1 U13531 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n11647) );
  INV_X1 U13532 ( .A(n13734), .ZN(n11645) );
  NAND2_X1 U13533 ( .A1(n11645), .A2(n11644), .ZN(n11646) );
  OAI21_X1 U13534 ( .B1(P3_U3897), .B2(n11647), .A(n11646), .ZN(P3_U3520) );
  NAND2_X1 U13535 ( .A1(n11648), .A2(n14040), .ZN(n16424) );
  NOR2_X1 U13536 ( .A1(n16424), .A2(n12920), .ZN(n11658) );
  INV_X1 U13537 ( .A(n11649), .ZN(n11650) );
  AOI21_X1 U13538 ( .B1(n12930), .B2(n11651), .A(n11650), .ZN(n11659) );
  OAI21_X1 U13539 ( .B1(n11653), .B2(n12930), .A(n11652), .ZN(n11656) );
  OAI22_X1 U13540 ( .A1(n11654), .A2(n13970), .B1(n11501), .B2(n13880), .ZN(
        n11655) );
  AOI21_X1 U13541 ( .B1(n11656), .B2(n13973), .A(n11655), .ZN(n11657) );
  OAI21_X1 U13542 ( .B1(n11659), .B2(n14015), .A(n11657), .ZN(n16425) );
  AOI211_X1 U13543 ( .C1(n13980), .C2(P3_REG3_REG_2__SCAN_IN), .A(n11658), .B(
        n16425), .ZN(n11661) );
  INV_X1 U13544 ( .A(n11659), .ZN(n16427) );
  AOI22_X1 U13545 ( .A1(n16427), .A2(n13846), .B1(n13910), .B2(
        P3_REG2_REG_2__SCAN_IN), .ZN(n11660) );
  OAI21_X1 U13546 ( .B1(n11661), .B2(n13958), .A(n11660), .ZN(P3_U3231) );
  INV_X1 U13547 ( .A(n11662), .ZN(n11663) );
  INV_X1 U13548 ( .A(n11720), .ZN(n11675) );
  NAND2_X1 U13549 ( .A1(P3_REG2_REG_9__SCAN_IN), .A2(n11664), .ZN(n11722) );
  OAI21_X1 U13550 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n11664), .A(n11722), .ZN(
        n11686) );
  OR2_X1 U13551 ( .A1(n11665), .A2(n12249), .ZN(n11666) );
  INV_X1 U13552 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n16542) );
  AOI21_X1 U13553 ( .B1(n11669), .B2(n16542), .A(n11726), .ZN(n11673) );
  INV_X1 U13554 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11670) );
  NOR2_X1 U13555 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11670), .ZN(n12464) );
  INV_X1 U13556 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n16257) );
  NOR2_X1 U13557 ( .A1(n16364), .A2(n16257), .ZN(n11671) );
  AOI211_X1 U13558 ( .C1(n13707), .C2(n11675), .A(n12464), .B(n11671), .ZN(
        n11672) );
  OAI21_X1 U13559 ( .B1(n11673), .B2(n16374), .A(n11672), .ZN(n11685) );
  MUX2_X1 U13560 ( .A(n11674), .B(n16542), .S(n7429), .Z(n11676) );
  NAND2_X1 U13561 ( .A1(n11676), .A2(n11675), .ZN(n11732) );
  INV_X1 U13562 ( .A(n11676), .ZN(n11677) );
  NAND2_X1 U13563 ( .A1(n11677), .A2(n11720), .ZN(n11678) );
  NAND2_X1 U13564 ( .A1(n11732), .A2(n11678), .ZN(n11679) );
  INV_X1 U13565 ( .A(n11740), .ZN(n11683) );
  NAND3_X1 U13566 ( .A1(n11681), .A2(n11680), .A3(n11679), .ZN(n11682) );
  AOI21_X1 U13567 ( .B1(n11683), .B2(n11682), .A(n16376), .ZN(n11684) );
  AOI211_X1 U13568 ( .C1(n13712), .C2(n11686), .A(n11685), .B(n11684), .ZN(
        n11687) );
  INV_X1 U13569 ( .A(n11687), .ZN(P3_U3191) );
  MUX2_X1 U13570 ( .A(n10951), .B(n11688), .S(n16587), .Z(n11692) );
  NAND2_X1 U13571 ( .A1(n16587), .A2(n16485), .ZN(n14063) );
  INV_X1 U13572 ( .A(n14063), .ZN(n16539) );
  AOI22_X1 U13573 ( .A1(n11690), .A2(n16539), .B1(n11689), .B2(n10089), .ZN(
        n11691) );
  NAND2_X1 U13574 ( .A1(n11692), .A2(n11691), .ZN(P3_U3463) );
  XOR2_X1 U13575 ( .A(n11694), .B(n11693), .Z(n11699) );
  INV_X1 U13576 ( .A(n12223), .ZN(n12082) );
  AOI22_X1 U13577 ( .A1(n14701), .A2(n14726), .B1(n14702), .B2(n14724), .ZN(
        n11697) );
  INV_X1 U13578 ( .A(n11695), .ZN(n12080) );
  AOI22_X1 U13579 ( .A1(n14700), .A2(n12080), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11696) );
  OAI211_X1 U13580 ( .C1(n12082), .C2(n14705), .A(n11697), .B(n11696), .ZN(
        n11698) );
  AOI21_X1 U13581 ( .B1(n11699), .B2(n14707), .A(n11698), .ZN(n11700) );
  INV_X1 U13582 ( .A(n11700), .ZN(P2_U3208) );
  INV_X1 U13583 ( .A(n13153), .ZN(n12728) );
  OAI222_X1 U13584 ( .A1(n15519), .A2(P1_U3086), .B1(n15990), .B2(n12728), 
        .C1(n11701), .C2(n15992), .ZN(P1_U3336) );
  INV_X1 U13585 ( .A(SI_23_), .ZN(n11705) );
  NAND2_X1 U13586 ( .A1(n11703), .A2(n11702), .ZN(n11704) );
  OAI211_X1 U13587 ( .C1(n11705), .C2(n14150), .A(n11704), .B(n12965), .ZN(
        P3_U3272) );
  INV_X1 U13588 ( .A(n11953), .ZN(n11717) );
  INV_X4 U13589 ( .A(n13425), .ZN(n13428) );
  XNOR2_X1 U13590 ( .A(n11706), .B(n13428), .ZN(n12155) );
  XNOR2_X1 U13591 ( .A(n12155), .B(n12163), .ZN(n11711) );
  INV_X1 U13592 ( .A(n11707), .ZN(n11708) );
  NAND2_X1 U13593 ( .A1(n11709), .A2(n11708), .ZN(n11710) );
  OAI21_X1 U13594 ( .B1(n11711), .B2(n11710), .A(n12157), .ZN(n11712) );
  NAND2_X1 U13595 ( .A1(n11712), .A2(n13576), .ZN(n11716) );
  OAI22_X1 U13596 ( .A1(n13582), .A2(n9997), .B1(n12384), .B2(n13593), .ZN(
        n11713) );
  AOI211_X1 U13597 ( .C1(n13589), .C2(n13485), .A(n11714), .B(n11713), .ZN(
        n11715) );
  OAI211_X1 U13598 ( .C1(n13448), .C2(n11717), .A(n11716), .B(n11715), .ZN(
        P3_U3167) );
  INV_X1 U13599 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11718) );
  MUX2_X1 U13600 ( .A(n11718), .B(P3_REG2_REG_10__SCAN_IN), .S(n11773), .Z(
        n11719) );
  INV_X1 U13601 ( .A(n11719), .ZN(n11725) );
  NAND2_X1 U13602 ( .A1(n11721), .A2(n11720), .ZN(n11723) );
  NAND2_X1 U13603 ( .A1(n11723), .A2(n11722), .ZN(n11724) );
  NAND2_X1 U13604 ( .A1(n11725), .A2(n11724), .ZN(n11774) );
  OAI21_X1 U13605 ( .B1(n11725), .B2(n11724), .A(n11774), .ZN(n11744) );
  NOR2_X1 U13606 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14272), .ZN(n12553) );
  NAND2_X1 U13607 ( .A1(n11773), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n11764) );
  OAI21_X1 U13608 ( .B1(n11773), .B2(P3_REG1_REG_10__SCAN_IN), .A(n11764), 
        .ZN(n11727) );
  AOI21_X1 U13609 ( .B1(n11728), .B2(n11727), .A(n11766), .ZN(n11729) );
  NOR2_X1 U13610 ( .A1(n16374), .A2(n11729), .ZN(n11730) );
  AOI211_X1 U13611 ( .C1(n16036), .C2(P3_ADDR_REG_10__SCAN_IN), .A(n12553), 
        .B(n11730), .ZN(n11731) );
  OAI21_X1 U13612 ( .B1(n11773), .B2(n16367), .A(n11731), .ZN(n11743) );
  INV_X1 U13613 ( .A(n11732), .ZN(n11739) );
  INV_X1 U13614 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11733) );
  MUX2_X1 U13615 ( .A(n11718), .B(n11733), .S(n7429), .Z(n11735) );
  INV_X1 U13616 ( .A(n11773), .ZN(n11734) );
  NAND2_X1 U13617 ( .A1(n11735), .A2(n11734), .ZN(n11768) );
  INV_X1 U13618 ( .A(n11735), .ZN(n11736) );
  NAND2_X1 U13619 ( .A1(n11736), .A2(n11773), .ZN(n11737) );
  AND2_X1 U13620 ( .A1(n11768), .A2(n11737), .ZN(n11738) );
  OR3_X1 U13621 ( .A1(n11740), .A2(n11739), .A3(n11738), .ZN(n11741) );
  AOI21_X1 U13622 ( .B1(n11769), .B2(n11741), .A(n16376), .ZN(n11742) );
  AOI211_X1 U13623 ( .C1(n13712), .C2(n11744), .A(n11743), .B(n11742), .ZN(
        n11745) );
  INV_X1 U13624 ( .A(n11745), .ZN(P3_U3192) );
  OR2_X1 U13625 ( .A1(n11746), .A2(n12812), .ZN(n11747) );
  NAND2_X1 U13626 ( .A1(n11748), .A2(n11747), .ZN(n12119) );
  NAND2_X1 U13627 ( .A1(n12119), .A2(n14052), .ZN(n11759) );
  NAND2_X1 U13628 ( .A1(n11947), .A2(n11750), .ZN(n11751) );
  NAND2_X1 U13629 ( .A1(n11751), .A2(n12812), .ZN(n11753) );
  NAND3_X1 U13630 ( .A1(n11753), .A2(n13973), .A3(n11752), .ZN(n11757) );
  OAI22_X1 U13631 ( .A1(n12388), .A2(n13880), .B1(n11754), .B2(n13970), .ZN(
        n11755) );
  INV_X1 U13632 ( .A(n11755), .ZN(n11756) );
  AND2_X1 U13633 ( .A1(n11757), .A2(n11756), .ZN(n11758) );
  NAND2_X1 U13634 ( .A1(n11759), .A2(n11758), .ZN(n12122) );
  INV_X1 U13635 ( .A(n12122), .ZN(n11763) );
  INV_X1 U13636 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n11760) );
  OAI22_X1 U13637 ( .A1(n14139), .A2(n12814), .B1(n16590), .B2(n11760), .ZN(
        n11761) );
  AOI21_X1 U13638 ( .B1(n12119), .B2(n14134), .A(n11761), .ZN(n11762) );
  OAI21_X1 U13639 ( .B1(n11763), .B2(n16588), .A(n11762), .ZN(P3_U3408) );
  INV_X1 U13640 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n16586) );
  INV_X1 U13641 ( .A(n11764), .ZN(n11765) );
  AOI21_X1 U13642 ( .B1(n16586), .B2(n11767), .A(n11887), .ZN(n11785) );
  NAND2_X1 U13643 ( .A1(n11769), .A2(n11768), .ZN(n11771) );
  MUX2_X1 U13644 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n7429), .Z(n11892) );
  XNOR2_X1 U13645 ( .A(n11892), .B(n11893), .ZN(n11770) );
  NAND2_X1 U13646 ( .A1(n11771), .A2(n11770), .ZN(n11899) );
  OAI21_X1 U13647 ( .B1(n11771), .B2(n11770), .A(n11899), .ZN(n11772) );
  NAND2_X1 U13648 ( .A1(n11772), .A2(n11900), .ZN(n11784) );
  NAND2_X1 U13649 ( .A1(n11773), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n11775) );
  NAND2_X1 U13650 ( .A1(n11775), .A2(n11774), .ZN(n11903) );
  XNOR2_X1 U13651 ( .A(n11903), .B(n11893), .ZN(n11776) );
  NAND2_X1 U13652 ( .A1(P3_REG2_REG_11__SCAN_IN), .A2(n11776), .ZN(n11905) );
  OAI21_X1 U13653 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n11776), .A(n11905), 
        .ZN(n11782) );
  INV_X1 U13654 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n11780) );
  NAND2_X1 U13655 ( .A1(n13707), .A2(n11893), .ZN(n11779) );
  INV_X1 U13656 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11777) );
  NOR2_X1 U13657 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11777), .ZN(n12662) );
  INV_X1 U13658 ( .A(n12662), .ZN(n11778) );
  OAI211_X1 U13659 ( .C1(n11780), .C2(n16364), .A(n11779), .B(n11778), .ZN(
        n11781) );
  AOI21_X1 U13660 ( .B1(n11782), .B2(n13712), .A(n11781), .ZN(n11783) );
  OAI211_X1 U13661 ( .C1(n11785), .C2(n16374), .A(n11784), .B(n11783), .ZN(
        P3_U3193) );
  INV_X1 U13662 ( .A(n16507), .ZN(n12075) );
  OR2_X1 U13663 ( .A1(n11787), .A2(n12075), .ZN(n11796) );
  NAND2_X1 U13664 ( .A1(n14829), .A2(n11796), .ZN(n16417) );
  OAI22_X1 U13665 ( .A1(n14926), .A2(n11788), .B1(n10708), .B2(n14922), .ZN(
        n11789) );
  AOI21_X1 U13666 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n14992), .A(n11789), .ZN(
        n11790) );
  OAI21_X1 U13667 ( .B1(n11791), .B2(n16515), .A(n11790), .ZN(n11792) );
  AOI21_X1 U13668 ( .B1(n11793), .B2(n16417), .A(n11792), .ZN(n11794) );
  OAI21_X1 U13669 ( .B1(n16522), .B2(n11795), .A(n11794), .ZN(P2_U3263) );
  INV_X1 U13670 ( .A(n13176), .ZN(n12046) );
  OAI222_X1 U13671 ( .A1(P1_U3086), .A2(n12993), .B1(n15990), .B2(n12046), 
        .C1(n13177), .C2(n15992), .ZN(P1_U3335) );
  MUX2_X1 U13672 ( .A(n10261), .B(n11797), .S(n14954), .Z(n11804) );
  INV_X1 U13673 ( .A(n11798), .ZN(n11800) );
  OAI22_X1 U13674 ( .A1(n14926), .A2(n11800), .B1(n11799), .B2(n14922), .ZN(
        n11801) );
  AOI21_X1 U13675 ( .B1(n16419), .B2(n11802), .A(n11801), .ZN(n11803) );
  OAI211_X1 U13676 ( .C1(n14892), .C2(n11805), .A(n11804), .B(n11803), .ZN(
        P2_U3260) );
  INV_X1 U13677 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11820) );
  INV_X1 U13678 ( .A(n11806), .ZN(n11807) );
  AOI21_X1 U13679 ( .B1(n11810), .B2(n11808), .A(n11807), .ZN(n16548) );
  OAI21_X1 U13680 ( .B1(n11811), .B2(n11810), .A(n11809), .ZN(n11814) );
  NOR2_X1 U13681 ( .A1(n16548), .A2(n16454), .ZN(n11812) );
  AOI211_X1 U13682 ( .C1(n16458), .C2(n11814), .A(n11813), .B(n11812), .ZN(
        n16553) );
  INV_X1 U13683 ( .A(n11815), .ZN(n11817) );
  AOI211_X1 U13684 ( .C1(n13078), .C2(n11817), .A(n15915), .B(n11816), .ZN(
        n16551) );
  AOI21_X1 U13685 ( .B1(n16490), .B2(n13078), .A(n16551), .ZN(n11818) );
  OAI211_X1 U13686 ( .C1(n16548), .C2(n16493), .A(n16553), .B(n11818), .ZN(
        n11821) );
  NAND2_X1 U13687 ( .A1(n11821), .A2(n16570), .ZN(n11819) );
  OAI21_X1 U13688 ( .B1(n16570), .B2(n11820), .A(n11819), .ZN(P1_U3486) );
  NAND2_X1 U13689 ( .A1(n11821), .A2(n16469), .ZN(n11822) );
  OAI21_X1 U13690 ( .B1(n16469), .B2(n11823), .A(n11822), .ZN(P1_U3537) );
  INV_X1 U13691 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11824) );
  XNOR2_X1 U13692 ( .A(n16102), .B(n11824), .ZN(n16103) );
  NAND2_X1 U13693 ( .A1(n11836), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n11828) );
  XNOR2_X1 U13694 ( .A(n16086), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n16093) );
  AOI21_X1 U13695 ( .B1(n11837), .B2(P2_REG1_REG_14__SCAN_IN), .A(n11825), 
        .ZN(n11826) );
  XOR2_X1 U13696 ( .A(n16079), .B(n11826), .Z(n16080) );
  INV_X1 U13697 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n11827) );
  OAI22_X1 U13698 ( .A1(n16080), .A2(n11827), .B1(n11826), .B2(n11842), .ZN(
        n16094) );
  NAND2_X1 U13699 ( .A1(n16093), .A2(n16094), .ZN(n16092) );
  NAND2_X1 U13700 ( .A1(n11828), .A2(n16092), .ZN(n16104) );
  AND2_X1 U13701 ( .A1(n16102), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n11829) );
  AOI21_X1 U13702 ( .B1(n16103), .B2(n16104), .A(n11829), .ZN(n11830) );
  XNOR2_X1 U13703 ( .A(n11830), .B(n16115), .ZN(n16116) );
  INV_X1 U13704 ( .A(n11830), .ZN(n11831) );
  AOI22_X1 U13705 ( .A1(n16116), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n16115), 
        .B2(n11831), .ZN(n11833) );
  XNOR2_X1 U13706 ( .A(n11851), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n11832) );
  XNOR2_X1 U13707 ( .A(n11833), .B(n11832), .ZN(n11859) );
  OR2_X1 U13708 ( .A1(n16102), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11834) );
  NAND2_X1 U13709 ( .A1(n16102), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11846) );
  AND2_X1 U13710 ( .A1(n11834), .A2(n11846), .ZN(n16101) );
  NAND2_X1 U13711 ( .A1(n11836), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11845) );
  NOR2_X1 U13712 ( .A1(n11836), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11835) );
  AOI21_X1 U13713 ( .B1(n11836), .B2(P2_REG2_REG_16__SCAN_IN), .A(n11835), 
        .ZN(n16090) );
  INV_X1 U13714 ( .A(n11838), .ZN(n11841) );
  OAI21_X1 U13715 ( .B1(n11838), .B2(P2_REG2_REG_14__SCAN_IN), .A(n11837), 
        .ZN(n11839) );
  OAI21_X1 U13716 ( .B1(n11841), .B2(n11840), .A(n11839), .ZN(n11843) );
  NAND2_X1 U13717 ( .A1(n16079), .A2(n11843), .ZN(n11844) );
  XNOR2_X1 U13718 ( .A(n11843), .B(n11842), .ZN(n16078) );
  NAND2_X1 U13719 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n16078), .ZN(n16077) );
  NAND2_X1 U13720 ( .A1(n11844), .A2(n16077), .ZN(n16091) );
  NAND2_X1 U13721 ( .A1(n16090), .A2(n16091), .ZN(n16089) );
  NAND2_X1 U13722 ( .A1(n11845), .A2(n16089), .ZN(n16100) );
  NAND2_X1 U13723 ( .A1(n16101), .A2(n16100), .ZN(n16099) );
  AND2_X1 U13724 ( .A1(n16099), .A2(n11846), .ZN(n11848) );
  NAND2_X1 U13725 ( .A1(n11848), .A2(n11847), .ZN(n11849) );
  OAI21_X1 U13726 ( .B1(n11848), .B2(n11847), .A(n11849), .ZN(n16112) );
  NOR2_X1 U13727 ( .A1(n16112), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n16111) );
  INV_X1 U13728 ( .A(n11849), .ZN(n11850) );
  NOR2_X1 U13729 ( .A1(n16111), .A2(n11850), .ZN(n11853) );
  MUX2_X1 U13730 ( .A(n8560), .B(P2_REG2_REG_19__SCAN_IN), .S(n11851), .Z(
        n11852) );
  XNOR2_X1 U13731 ( .A(n11853), .B(n11852), .ZN(n11856) );
  AND2_X1 U13732 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14184) );
  AOI21_X1 U13733 ( .B1(n16110), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n14184), 
        .ZN(n11854) );
  OAI21_X1 U13734 ( .B1(n16127), .B2(n12727), .A(n11854), .ZN(n11855) );
  AOI21_X1 U13735 ( .B1(n16152), .B2(n11856), .A(n11855), .ZN(n11857) );
  OAI21_X1 U13736 ( .B1(n11859), .B2(n11858), .A(n11857), .ZN(P2_U3233) );
  INV_X1 U13737 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11883) );
  OR2_X1 U13738 ( .A1(n13082), .A2(n15375), .ZN(n11860) );
  NAND2_X1 U13739 ( .A1(n11862), .A2(n13289), .ZN(n11865) );
  AOI22_X1 U13740 ( .A1(n11863), .A2(n13154), .B1(n13155), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n11864) );
  XNOR2_X1 U13741 ( .A(n13086), .B(n15374), .ZN(n13324) );
  NAND2_X1 U13742 ( .A1(n11866), .A2(n13324), .ZN(n11867) );
  NAND2_X1 U13743 ( .A1(n11958), .A2(n11867), .ZN(n16598) );
  NOR2_X1 U13744 ( .A1(n13324), .A2(n7564), .ZN(n11869) );
  AOI21_X1 U13745 ( .B1(n11870), .B2(n11869), .A(n16558), .ZN(n11880) );
  NAND2_X1 U13746 ( .A1(n13170), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n11877) );
  OR2_X1 U13747 ( .A1(n13256), .A2(n10835), .ZN(n11876) );
  NAND2_X1 U13748 ( .A1(n11871), .A2(n12183), .ZN(n11872) );
  NAND2_X1 U13749 ( .A1(n11969), .A2(n11872), .ZN(n12182) );
  OR2_X1 U13750 ( .A1(n13282), .A2(n12182), .ZN(n11875) );
  INV_X1 U13751 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11873) );
  OR2_X1 U13752 ( .A1(n13284), .A2(n11873), .ZN(n11874) );
  NAND4_X1 U13753 ( .A1(n11877), .A2(n11876), .A3(n11875), .A4(n11874), .ZN(
        n15373) );
  NAND2_X1 U13754 ( .A1(n15789), .A2(n15373), .ZN(n11879) );
  NAND2_X1 U13755 ( .A1(n15787), .A2(n15375), .ZN(n11878) );
  NAND2_X1 U13756 ( .A1(n11879), .A2(n11878), .ZN(n12060) );
  AOI21_X1 U13757 ( .B1(n11966), .B2(n11880), .A(n12060), .ZN(n16604) );
  INV_X1 U13758 ( .A(n11981), .ZN(n11983) );
  AOI211_X1 U13759 ( .C1(n13086), .C2(n7563), .A(n15915), .B(n11983), .ZN(
        n16602) );
  AOI21_X1 U13760 ( .B1(n16490), .B2(n13086), .A(n16602), .ZN(n11881) );
  OAI211_X1 U13761 ( .C1(n16435), .C2(n16598), .A(n16604), .B(n11881), .ZN(
        n11884) );
  NAND2_X1 U13762 ( .A1(n11884), .A2(n16570), .ZN(n11882) );
  OAI21_X1 U13763 ( .B1(n16570), .B2(n11883), .A(n11882), .ZN(P1_U3492) );
  NAND2_X1 U13764 ( .A1(n11884), .A2(n16469), .ZN(n11885) );
  OAI21_X1 U13765 ( .B1(n16469), .B2(n11600), .A(n11885), .ZN(P1_U3539) );
  OR2_X1 U13766 ( .A1(n11895), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n11888) );
  NAND2_X1 U13767 ( .A1(n11895), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12441) );
  AND2_X1 U13768 ( .A1(n11888), .A2(n12441), .ZN(n11897) );
  INV_X1 U13769 ( .A(n11897), .ZN(n11890) );
  INV_X1 U13770 ( .A(n12435), .ZN(n11889) );
  AOI21_X1 U13771 ( .B1(n11891), .B2(n11890), .A(n11889), .ZN(n11917) );
  INV_X1 U13772 ( .A(n11892), .ZN(n11894) );
  NAND2_X1 U13773 ( .A1(n11894), .A2(n11893), .ZN(n11898) );
  AND2_X1 U13774 ( .A1(n11899), .A2(n11898), .ZN(n11902) );
  INV_X1 U13775 ( .A(n11895), .ZN(n11909) );
  INV_X1 U13776 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n13978) );
  NAND2_X1 U13777 ( .A1(n11895), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12442) );
  INV_X1 U13778 ( .A(n12442), .ZN(n11896) );
  AOI21_X1 U13779 ( .B1(n11909), .B2(n13978), .A(n11896), .ZN(n11908) );
  MUX2_X1 U13780 ( .A(n11908), .B(n11897), .S(n7429), .Z(n11901) );
  NAND3_X1 U13781 ( .A1(n11899), .A2(n11898), .A3(n11901), .ZN(n12444) );
  OAI211_X1 U13782 ( .C1(n11902), .C2(n11901), .A(n11900), .B(n12444), .ZN(
        n11916) );
  NAND2_X1 U13783 ( .A1(n11904), .A2(n11903), .ZN(n11906) );
  NAND2_X1 U13784 ( .A1(n11906), .A2(n11905), .ZN(n11907) );
  OAI21_X1 U13785 ( .B1(n11908), .B2(n11907), .A(n12438), .ZN(n11914) );
  INV_X1 U13786 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n11912) );
  NAND2_X1 U13787 ( .A1(n13707), .A2(n11909), .ZN(n11911) );
  INV_X1 U13788 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11910) );
  OR2_X1 U13789 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11910), .ZN(n12621) );
  OAI211_X1 U13790 ( .C1(n11912), .C2(n16364), .A(n11911), .B(n12621), .ZN(
        n11913) );
  AOI21_X1 U13791 ( .B1(n11914), .B2(n13712), .A(n11913), .ZN(n11915) );
  OAI211_X1 U13792 ( .C1(n11917), .C2(n16374), .A(n11916), .B(n11915), .ZN(
        P3_U3194) );
  XNOR2_X1 U13793 ( .A(n11919), .B(n11918), .ZN(n16502) );
  INV_X1 U13794 ( .A(n16502), .ZN(n11937) );
  INV_X1 U13795 ( .A(n11920), .ZN(n11921) );
  AOI21_X1 U13796 ( .B1(n11923), .B2(n11922), .A(n11921), .ZN(n11926) );
  AOI22_X1 U13797 ( .A1(n14913), .A2(n14729), .B1(n14731), .B2(n14911), .ZN(
        n11925) );
  NAND2_X1 U13798 ( .A1(n16502), .A2(n16507), .ZN(n11924) );
  OAI211_X1 U13799 ( .C1(n11926), .C2(n14949), .A(n11925), .B(n11924), .ZN(
        n16500) );
  NAND2_X1 U13800 ( .A1(n16500), .A2(n14954), .ZN(n11936) );
  OAI21_X1 U13801 ( .B1(n11927), .B2(n16499), .A(n14930), .ZN(n11929) );
  OR2_X1 U13802 ( .A1(n11929), .A2(n11928), .ZN(n16498) );
  NOR2_X1 U13803 ( .A1(n14926), .A2(n16498), .ZN(n11933) );
  OAI22_X1 U13804 ( .A1(n14954), .A2(n11931), .B1(n11930), .B2(n14922), .ZN(
        n11932) );
  AOI211_X1 U13805 ( .C1(n16419), .C2(n11934), .A(n11933), .B(n11932), .ZN(
        n11935) );
  OAI211_X1 U13806 ( .C1(n11937), .C2(n14829), .A(n11936), .B(n11935), .ZN(
        P2_U3259) );
  OR2_X1 U13807 ( .A1(n11938), .A2(n12925), .ZN(n11939) );
  NAND2_X1 U13808 ( .A1(n11940), .A2(n11939), .ZN(n16484) );
  INV_X1 U13809 ( .A(n16484), .ZN(n11956) );
  NAND2_X1 U13810 ( .A1(n16484), .A2(n14052), .ZN(n11951) );
  NAND2_X1 U13811 ( .A1(n11942), .A2(n11941), .ZN(n11944) );
  AND2_X1 U13812 ( .A1(n11944), .A2(n11943), .ZN(n11945) );
  NAND2_X1 U13813 ( .A1(n11945), .A2(n12925), .ZN(n11946) );
  NAND2_X1 U13814 ( .A1(n11947), .A2(n11946), .ZN(n11948) );
  NAND2_X1 U13815 ( .A1(n11948), .A2(n13973), .ZN(n11950) );
  AOI22_X1 U13816 ( .A1(n13485), .A2(n13954), .B1(n13967), .B2(n13605), .ZN(
        n11949) );
  NAND3_X1 U13817 ( .A1(n11951), .A2(n11950), .A3(n11949), .ZN(n16482) );
  MUX2_X1 U13818 ( .A(n16482), .B(P3_REG2_REG_5__SCAN_IN), .S(n13910), .Z(
        n11952) );
  INV_X1 U13819 ( .A(n11952), .ZN(n11955) );
  AOI22_X1 U13820 ( .A1(n13981), .A2(n11706), .B1(n11953), .B2(n13980), .ZN(
        n11954) );
  OAI211_X1 U13821 ( .C1(n11956), .C2(n13984), .A(n11955), .B(n11954), .ZN(
        P3_U3228) );
  NAND2_X1 U13822 ( .A1(n13086), .A2(n15374), .ZN(n11957) );
  AND2_X2 U13823 ( .A1(n11958), .A2(n11957), .ZN(n11964) );
  NAND2_X1 U13824 ( .A1(n11959), .A2(n13289), .ZN(n11962) );
  AOI22_X1 U13825 ( .A1(n13155), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n13154), 
        .B2(n11960), .ZN(n11961) );
  XNOR2_X1 U13826 ( .A(n13090), .B(n15373), .ZN(n13326) );
  INV_X1 U13827 ( .A(n13326), .ZN(n11963) );
  OAI21_X1 U13828 ( .B1(n11964), .B2(n11963), .A(n12020), .ZN(n12234) );
  INV_X1 U13829 ( .A(n12234), .ZN(n11988) );
  OR2_X1 U13830 ( .A1(n13086), .A2(n12050), .ZN(n11965) );
  NAND2_X1 U13831 ( .A1(n11966), .A2(n11965), .ZN(n11967) );
  NAND2_X1 U13832 ( .A1(n11967), .A2(n13326), .ZN(n11998) );
  OAI211_X1 U13833 ( .C1(n11967), .C2(n13326), .A(n11998), .B(n16458), .ZN(
        n11980) );
  INV_X1 U13834 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n11968) );
  NAND2_X1 U13835 ( .A1(n11969), .A2(n11968), .ZN(n11970) );
  NAND2_X1 U13836 ( .A1(n12008), .A2(n11970), .ZN(n12363) );
  OR2_X1 U13837 ( .A1(n13282), .A2(n12363), .ZN(n11977) );
  INV_X1 U13838 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11971) );
  OR2_X1 U13839 ( .A1(n13279), .A2(n11971), .ZN(n11976) );
  INV_X1 U13840 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11972) );
  OR2_X1 U13841 ( .A1(n13256), .A2(n11972), .ZN(n11975) );
  OR2_X1 U13842 ( .A1(n13284), .A2(n11973), .ZN(n11974) );
  NAND4_X1 U13843 ( .A1(n11977), .A2(n11976), .A3(n11975), .A4(n11974), .ZN(
        n15372) );
  NAND2_X1 U13844 ( .A1(n15789), .A2(n15372), .ZN(n11979) );
  NAND2_X1 U13845 ( .A1(n15787), .A2(n15374), .ZN(n11978) );
  AND2_X1 U13846 ( .A1(n11979), .A2(n11978), .ZN(n12184) );
  NAND2_X1 U13847 ( .A1(n11980), .A2(n12184), .ZN(n12232) );
  NAND2_X1 U13848 ( .A1(n12232), .A2(n15812), .ZN(n11987) );
  OAI22_X1 U13849 ( .A1(n15812), .A2(n10835), .B1(n12182), .B2(n16395), .ZN(
        n11985) );
  INV_X1 U13850 ( .A(n13090), .ZN(n12231) );
  INV_X1 U13851 ( .A(n12005), .ZN(n11982) );
  OAI211_X1 U13852 ( .C1(n12231), .C2(n11983), .A(n11982), .B(n15910), .ZN(
        n12230) );
  NOR2_X1 U13853 ( .A1(n12230), .A2(n15780), .ZN(n11984) );
  AOI211_X1 U13854 ( .C1(n16525), .C2(n13090), .A(n11985), .B(n11984), .ZN(
        n11986) );
  OAI211_X1 U13855 ( .C1(n16597), .C2(n11988), .A(n11987), .B(n11986), .ZN(
        P1_U3281) );
  OAI22_X1 U13856 ( .A1(n14926), .A2(n11989), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14922), .ZN(n11992) );
  NOR2_X1 U13857 ( .A1(n16515), .A2(n11990), .ZN(n11991) );
  AOI211_X1 U13858 ( .C1(n14992), .C2(P2_REG2_REG_3__SCAN_IN), .A(n11992), .B(
        n11991), .ZN(n11995) );
  NAND2_X1 U13859 ( .A1(n16417), .A2(n11993), .ZN(n11994) );
  OAI211_X1 U13860 ( .C1(n16522), .C2(n11996), .A(n11995), .B(n11994), .ZN(
        P2_U3262) );
  INV_X1 U13861 ( .A(n15373), .ZN(n12178) );
  OR2_X1 U13862 ( .A1(n13090), .A2(n12178), .ZN(n11997) );
  NAND2_X1 U13863 ( .A1(n11998), .A2(n11997), .ZN(n12004) );
  NAND2_X1 U13864 ( .A1(n11999), .A2(n13289), .ZN(n12002) );
  AOI22_X1 U13865 ( .A1(n13155), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n12000), 
        .B2(n13154), .ZN(n12001) );
  INV_X1 U13866 ( .A(n15372), .ZN(n12359) );
  XNOR2_X1 U13867 ( .A(n15940), .B(n12359), .ZN(n13328) );
  INV_X1 U13868 ( .A(n13328), .ZN(n12003) );
  OAI21_X1 U13869 ( .B1(n12004), .B2(n12003), .A(n12311), .ZN(n15944) );
  INV_X1 U13870 ( .A(n15940), .ZN(n12368) );
  OAI21_X1 U13871 ( .B1(n12005), .B2(n12368), .A(n15910), .ZN(n12006) );
  AND2_X2 U13872 ( .A1(n12005), .A2(n12368), .ZN(n12320) );
  NOR2_X1 U13873 ( .A1(n12006), .A2(n12320), .ZN(n15938) );
  INV_X1 U13874 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n12007) );
  AND2_X1 U13875 ( .A1(n12008), .A2(n12007), .ZN(n12009) );
  OR2_X1 U13876 ( .A1(n12009), .A2(n12321), .ZN(n12521) );
  OR2_X1 U13877 ( .A1(n13256), .A2(n11446), .ZN(n12012) );
  INV_X1 U13878 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n12010) );
  OR2_X1 U13879 ( .A1(n13284), .A2(n12010), .ZN(n12011) );
  AND2_X1 U13880 ( .A1(n12012), .A2(n12011), .ZN(n12014) );
  NAND2_X1 U13881 ( .A1(n13170), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n12013) );
  OAI211_X1 U13882 ( .C1(n13282), .C2(n12521), .A(n12014), .B(n12013), .ZN(
        n15371) );
  INV_X1 U13883 ( .A(n15371), .ZN(n15358) );
  OAI22_X1 U13884 ( .A1(n15358), .A2(n16389), .B1(n12178), .B2(n15805), .ZN(
        n15939) );
  INV_X1 U13885 ( .A(n12363), .ZN(n12015) );
  AOI22_X1 U13886 ( .A1(n15812), .A2(n15939), .B1(n12015), .B2(n16592), .ZN(
        n12017) );
  NAND2_X1 U13887 ( .A1(n16605), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n12016) );
  OAI211_X1 U13888 ( .C1(n12368), .C2(n16595), .A(n12017), .B(n12016), .ZN(
        n12018) );
  AOI21_X1 U13889 ( .B1(n15938), .B2(n16601), .A(n12018), .ZN(n12023) );
  OR2_X1 U13890 ( .A1(n13090), .A2(n15373), .ZN(n12019) );
  OAI21_X1 U13891 ( .B1(n12021), .B2(n13328), .A(n12317), .ZN(n15941) );
  NAND2_X1 U13892 ( .A1(n15941), .A2(n15818), .ZN(n12022) );
  OAI211_X1 U13893 ( .C1(n15944), .C2(n15821), .A(n12023), .B(n12022), .ZN(
        P1_U3280) );
  INV_X1 U13894 ( .A(n12033), .ZN(n12025) );
  NAND3_X1 U13895 ( .A1(n11549), .A2(n12025), .A3(n12024), .ZN(n12026) );
  AND2_X1 U13896 ( .A1(n12027), .A2(n12026), .ZN(n12028) );
  OAI222_X1 U13897 ( .A1(n14953), .A2(n12065), .B1(n14951), .B2(n12029), .C1(
        n14949), .C2(n12028), .ZN(n16534) );
  INV_X1 U13898 ( .A(n16534), .ZN(n12044) );
  INV_X1 U13899 ( .A(n12030), .ZN(n12031) );
  AOI21_X1 U13900 ( .B1(n12033), .B2(n12032), .A(n12031), .ZN(n16536) );
  AOI21_X1 U13901 ( .B1(n12035), .B2(n12034), .A(n14986), .ZN(n12037) );
  NAND2_X1 U13902 ( .A1(n12037), .A2(n12036), .ZN(n16533) );
  NOR2_X1 U13903 ( .A1(n16533), .A2(n14926), .ZN(n12042) );
  INV_X1 U13904 ( .A(n12038), .ZN(n12039) );
  AOI22_X1 U13905 ( .A1(n14992), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n12039), 
        .B2(n16511), .ZN(n12040) );
  OAI21_X1 U13906 ( .B1(n16515), .B2(n7947), .A(n12040), .ZN(n12041) );
  AOI211_X1 U13907 ( .C1(n16536), .C2(n16417), .A(n12042), .B(n12041), .ZN(
        n12043) );
  OAI21_X1 U13908 ( .B1(n12044), .B2(n14992), .A(n12043), .ZN(P2_U3257) );
  OAI222_X1 U13909 ( .A1(n15131), .A2(n12046), .B1(P2_U3088), .B2(n9155), .C1(
        n12045), .C2(n15133), .ZN(P2_U3307) );
  INV_X1 U13910 ( .A(n13086), .ZN(n16596) );
  NAND2_X1 U13911 ( .A1(n13086), .A2(n15255), .ZN(n12048) );
  NAND2_X1 U13912 ( .A1(n15374), .A2(n7432), .ZN(n12047) );
  NAND2_X1 U13913 ( .A1(n12048), .A2(n12047), .ZN(n12049) );
  XNOR2_X1 U13914 ( .A(n12049), .B(n15253), .ZN(n12170) );
  NOR2_X1 U13915 ( .A1(n12050), .A2(n15223), .ZN(n12051) );
  AOI21_X1 U13916 ( .B1(n13086), .B2(n7432), .A(n12051), .ZN(n12171) );
  XNOR2_X1 U13917 ( .A(n12170), .B(n12171), .ZN(n12056) );
  OR2_X1 U13918 ( .A1(n12053), .A2(n12052), .ZN(n12054) );
  OAI21_X1 U13919 ( .B1(n12056), .B2(n7556), .A(n12174), .ZN(n12057) );
  NAND2_X1 U13920 ( .A1(n12057), .A2(n15332), .ZN(n12062) );
  NOR2_X1 U13921 ( .A1(n15360), .A2(n16591), .ZN(n12058) );
  AOI211_X1 U13922 ( .C1(n15277), .C2(n12060), .A(n12059), .B(n12058), .ZN(
        n12061) );
  OAI211_X1 U13923 ( .C1(n16596), .C2(n15340), .A(n12062), .B(n12061), .ZN(
        P1_U3236) );
  OR2_X1 U13924 ( .A1(n12095), .A2(n12065), .ZN(n12063) );
  NAND2_X1 U13925 ( .A1(n12064), .A2(n12063), .ZN(n12067) );
  NAND2_X1 U13926 ( .A1(n12095), .A2(n12065), .ZN(n12066) );
  NAND2_X1 U13927 ( .A1(n12067), .A2(n12066), .ZN(n12142) );
  INV_X1 U13928 ( .A(n12073), .ZN(n12068) );
  OAI21_X1 U13929 ( .B1(n7567), .B2(n12068), .A(n12192), .ZN(n12077) );
  OR2_X1 U13930 ( .A1(n12151), .A2(n14726), .ZN(n12071) );
  OAI21_X1 U13931 ( .B1(n7558), .B2(n12073), .A(n12190), .ZN(n12226) );
  AOI22_X1 U13932 ( .A1(n14911), .A2(n14726), .B1(n14724), .B2(n14913), .ZN(
        n12074) );
  OAI21_X1 U13933 ( .B1(n12226), .B2(n12075), .A(n12074), .ZN(n12076) );
  AOI21_X1 U13934 ( .B1(n14981), .B2(n12077), .A(n12076), .ZN(n12225) );
  INV_X1 U13935 ( .A(n12078), .ZN(n12146) );
  INV_X1 U13936 ( .A(n12201), .ZN(n12079) );
  AOI211_X1 U13937 ( .C1(n12223), .C2(n12146), .A(n14873), .B(n12079), .ZN(
        n12222) );
  AOI22_X1 U13938 ( .A1(n14992), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n12080), 
        .B2(n16511), .ZN(n12081) );
  OAI21_X1 U13939 ( .B1(n12082), .B2(n16515), .A(n12081), .ZN(n12084) );
  NOR2_X1 U13940 ( .A1(n12226), .A2(n14829), .ZN(n12083) );
  AOI211_X1 U13941 ( .C1(n12222), .C2(n16508), .A(n12084), .B(n12083), .ZN(
        n12085) );
  OAI21_X1 U13942 ( .B1(n16522), .B2(n12225), .A(n12085), .ZN(P2_U3254) );
  NAND3_X1 U13943 ( .A1(n14629), .A2(n14671), .A3(n14724), .ZN(n12086) );
  OAI21_X1 U13944 ( .B1(n12087), .B2(n14686), .A(n12086), .ZN(n12089) );
  NAND2_X1 U13945 ( .A1(n12089), .A2(n12088), .ZN(n12094) );
  AOI22_X1 U13946 ( .A1(n14702), .A2(n14722), .B1(n14701), .B2(n14724), .ZN(
        n12091) );
  OAI211_X1 U13947 ( .C1(n12274), .C2(n14683), .A(n12091), .B(n12090), .ZN(
        n12092) );
  AOI21_X1 U13948 ( .B1(n12427), .B2(n14691), .A(n12092), .ZN(n12093) );
  OAI211_X1 U13949 ( .C1(n12135), .C2(n14686), .A(n12094), .B(n12093), .ZN(
        P2_U3206) );
  INV_X1 U13950 ( .A(n12095), .ZN(n12096) );
  NOR2_X1 U13951 ( .A1(n16515), .A2(n12096), .ZN(n12100) );
  OAI22_X1 U13952 ( .A1(n14954), .A2(n12098), .B1(n12097), .B2(n14922), .ZN(
        n12099) );
  AOI211_X1 U13953 ( .C1(n12101), .C2(n16508), .A(n12100), .B(n12099), .ZN(
        n12104) );
  NAND2_X1 U13954 ( .A1(n12102), .A2(n16519), .ZN(n12103) );
  OAI211_X1 U13955 ( .C1(n12105), .C2(n16522), .A(n12104), .B(n12103), .ZN(
        P2_U3256) );
  XNOR2_X1 U13956 ( .A(n12106), .B(n12924), .ZN(n12283) );
  NAND2_X1 U13957 ( .A1(n12283), .A2(n14052), .ZN(n12114) );
  XNOR2_X1 U13958 ( .A(n12108), .B(n12924), .ZN(n12112) );
  NAND2_X1 U13959 ( .A1(n13604), .A2(n13967), .ZN(n12110) );
  NAND2_X1 U13960 ( .A1(n13605), .A2(n13954), .ZN(n12109) );
  NAND2_X1 U13961 ( .A1(n12110), .A2(n12109), .ZN(n12111) );
  AOI21_X1 U13962 ( .B1(n12112), .B2(n13973), .A(n12111), .ZN(n12113) );
  AND2_X1 U13963 ( .A1(n12114), .A2(n12113), .ZN(n12284) );
  OAI22_X1 U13964 ( .A1(n14139), .A2(n12116), .B1(n16590), .B2(n12115), .ZN(
        n12117) );
  AOI21_X1 U13965 ( .B1(n12283), .B2(n14134), .A(n12117), .ZN(n12118) );
  OAI21_X1 U13966 ( .B1(n12284), .B2(n16588), .A(n12118), .ZN(P3_U3411) );
  MUX2_X1 U13967 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n12122), .S(n16587), .Z(
        n12121) );
  INV_X1 U13968 ( .A(n12119), .ZN(n12126) );
  OAI22_X1 U13969 ( .A1(n12126), .A2(n14063), .B1(n12814), .B2(n14051), .ZN(
        n12120) );
  OR2_X1 U13970 ( .A1(n12121), .A2(n12120), .ZN(P3_U3465) );
  MUX2_X1 U13971 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n12122), .S(n13977), .Z(
        n12123) );
  INV_X1 U13972 ( .A(n12123), .ZN(n12125) );
  AOI22_X1 U13973 ( .A1(n13981), .A2(n12164), .B1(n13980), .B2(n12161), .ZN(
        n12124) );
  OAI211_X1 U13974 ( .C1(n12126), .C2(n13984), .A(n12125), .B(n12124), .ZN(
        P3_U3227) );
  NAND2_X1 U13975 ( .A1(n14721), .A2(n14913), .ZN(n12128) );
  NAND2_X1 U13976 ( .A1(n14723), .A2(n14911), .ZN(n12127) );
  AND2_X1 U13977 ( .A1(n12128), .A2(n12127), .ZN(n12372) );
  OAI22_X1 U13978 ( .A1(n14650), .A2(n12372), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12129), .ZN(n12131) );
  INV_X1 U13979 ( .A(n12566), .ZN(n16617) );
  NOR2_X1 U13980 ( .A1(n16617), .A2(n14705), .ZN(n12130) );
  AOI211_X1 U13981 ( .C1(n14700), .C2(n12378), .A(n12131), .B(n12130), .ZN(
        n12137) );
  OAI22_X1 U13982 ( .A1(n12133), .A2(n14686), .B1(n12369), .B2(n14694), .ZN(
        n12134) );
  NAND3_X1 U13983 ( .A1(n12135), .A2(n8027), .A3(n12134), .ZN(n12136) );
  OAI211_X1 U13984 ( .C1(n12138), .C2(n14686), .A(n12137), .B(n12136), .ZN(
        P2_U3187) );
  INV_X1 U13985 ( .A(n13182), .ZN(n12140) );
  OAI222_X1 U13986 ( .A1(n12999), .A2(P1_U3086), .B1(n15990), .B2(n12140), 
        .C1(n13183), .C2(n15987), .ZN(P1_U3334) );
  OAI222_X1 U13987 ( .A1(n15133), .A2(n12141), .B1(n15123), .B2(n12140), .C1(
        P2_U3088), .C2(n12139), .ZN(P2_U3306) );
  XNOR2_X1 U13988 ( .A(n12142), .B(n12144), .ZN(n12143) );
  AOI222_X1 U13989 ( .A1(n14981), .A2(n12143), .B1(n14725), .B2(n14913), .C1(
        n14727), .C2(n14911), .ZN(n16572) );
  XNOR2_X1 U13990 ( .A(n12145), .B(n12144), .ZN(n16575) );
  OAI211_X1 U13991 ( .C1(n16573), .C2(n12147), .A(n12146), .B(n14930), .ZN(
        n16571) );
  OAI22_X1 U13992 ( .A1(n14954), .A2(n12149), .B1(n12148), .B2(n14922), .ZN(
        n12150) );
  AOI21_X1 U13993 ( .B1(n16419), .B2(n12151), .A(n12150), .ZN(n12152) );
  OAI21_X1 U13994 ( .B1(n16571), .B2(n14926), .A(n12152), .ZN(n12153) );
  AOI21_X1 U13995 ( .B1(n16575), .B2(n16417), .A(n12153), .ZN(n12154) );
  OAI21_X1 U13996 ( .B1(n16572), .B2(n14992), .A(n12154), .ZN(P2_U3255) );
  XNOR2_X1 U13997 ( .A(n12814), .B(n13428), .ZN(n12385) );
  XNOR2_X1 U13998 ( .A(n12385), .B(n13605), .ZN(n12160) );
  NAND2_X1 U13999 ( .A1(n12155), .A2(n11754), .ZN(n12156) );
  INV_X1 U14000 ( .A(n12387), .ZN(n12158) );
  AOI211_X1 U14001 ( .C1(n12160), .C2(n12159), .A(n13599), .B(n12158), .ZN(
        n12169) );
  INV_X1 U14002 ( .A(n12161), .ZN(n12167) );
  AOI21_X1 U14003 ( .B1(n12163), .B2(n13589), .A(n12162), .ZN(n12166) );
  AOI22_X1 U14004 ( .A1(n12394), .A2(n13566), .B1(n13596), .B2(n12164), .ZN(
        n12165) );
  OAI211_X1 U14005 ( .C1(n12167), .C2(n13448), .A(n12166), .B(n12165), .ZN(
        n12168) );
  OR2_X1 U14006 ( .A1(n12169), .A2(n12168), .ZN(P3_U3179) );
  INV_X1 U14007 ( .A(n12170), .ZN(n12172) );
  NAND2_X1 U14008 ( .A1(n12172), .A2(n12171), .ZN(n12173) );
  NAND2_X1 U14009 ( .A1(n13090), .A2(n15255), .ZN(n12176) );
  NAND2_X1 U14010 ( .A1(n15373), .A2(n7432), .ZN(n12175) );
  NAND2_X1 U14011 ( .A1(n12176), .A2(n12175), .ZN(n12177) );
  XNOR2_X1 U14012 ( .A(n12177), .B(n15253), .ZN(n12351) );
  NOR2_X1 U14013 ( .A1(n12178), .A2(n15223), .ZN(n12179) );
  AOI21_X1 U14014 ( .B1(n13090), .B2(n7432), .A(n12179), .ZN(n12352) );
  XNOR2_X1 U14015 ( .A(n12351), .B(n12352), .ZN(n12180) );
  OAI211_X1 U14016 ( .C1(n12181), .C2(n12180), .A(n12355), .B(n15332), .ZN(
        n12188) );
  INV_X1 U14017 ( .A(n12182), .ZN(n12186) );
  OAI22_X1 U14018 ( .A1(n15264), .A2(n12184), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12183), .ZN(n12185) );
  AOI21_X1 U14019 ( .B1(n12186), .B2(n15312), .A(n12185), .ZN(n12187) );
  OAI211_X1 U14020 ( .C1(n12231), .C2(n15340), .A(n12188), .B(n12187), .ZN(
        P1_U3224) );
  NAND2_X1 U14021 ( .A1(n12223), .A2(n14725), .ZN(n12189) );
  XNOR2_X1 U14022 ( .A(n12262), .B(n12194), .ZN(n16611) );
  NAND2_X1 U14023 ( .A1(n16611), .A2(n16507), .ZN(n12200) );
  OAI21_X1 U14024 ( .B1(n12194), .B2(n12193), .A(n12266), .ZN(n12198) );
  NAND2_X1 U14025 ( .A1(n14725), .A2(n14911), .ZN(n12196) );
  NAND2_X1 U14026 ( .A1(n14723), .A2(n14913), .ZN(n12195) );
  NAND2_X1 U14027 ( .A1(n12196), .A2(n12195), .ZN(n12197) );
  AOI21_X1 U14028 ( .B1(n12198), .B2(n14981), .A(n12197), .ZN(n12199) );
  AND2_X1 U14029 ( .A1(n12200), .A2(n12199), .ZN(n16613) );
  AOI21_X1 U14030 ( .B1(n12201), .B2(n16606), .A(n14986), .ZN(n12202) );
  NAND2_X1 U14031 ( .A1(n12202), .A2(n12273), .ZN(n16607) );
  OAI22_X1 U14032 ( .A1(n14954), .A2(n12203), .B1(n14631), .B2(n14922), .ZN(
        n12204) );
  AOI21_X1 U14033 ( .B1(n16419), .B2(n16606), .A(n12204), .ZN(n12205) );
  OAI21_X1 U14034 ( .B1(n16607), .B2(n14926), .A(n12205), .ZN(n12206) );
  AOI21_X1 U14035 ( .B1(n16611), .B2(n16519), .A(n12206), .ZN(n12207) );
  OAI21_X1 U14036 ( .B1(n16613), .B2(n16522), .A(n12207), .ZN(P2_U3253) );
  INV_X1 U14037 ( .A(n12208), .ZN(n12210) );
  NAND2_X1 U14038 ( .A1(n12210), .A2(n12209), .ZN(n12334) );
  OR2_X1 U14039 ( .A1(n13110), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n12211) );
  NAND2_X1 U14040 ( .A1(n13110), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n12336) );
  NAND2_X1 U14041 ( .A1(n12211), .A2(n12336), .ZN(n12333) );
  XNOR2_X1 U14042 ( .A(n12334), .B(n12333), .ZN(n12221) );
  NAND2_X1 U14043 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n15289)
         );
  XOR2_X1 U14044 ( .A(n13110), .B(P1_REG1_REG_16__SCAN_IN), .Z(n12216) );
  INV_X1 U14045 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n12325) );
  NAND2_X1 U14046 ( .A1(n12216), .A2(n12215), .ZN(n12339) );
  OAI211_X1 U14047 ( .C1(n12216), .C2(n12215), .A(n15517), .B(n12339), .ZN(
        n12217) );
  NAND2_X1 U14048 ( .A1(n15289), .A2(n12217), .ZN(n12219) );
  NOR2_X1 U14049 ( .A1(n15511), .A2(n12340), .ZN(n12218) );
  AOI211_X1 U14050 ( .C1(n16162), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n12219), 
        .B(n12218), .ZN(n12220) );
  OAI21_X1 U14051 ( .B1(n12221), .B2(n15512), .A(n12220), .ZN(P1_U3259) );
  AOI21_X1 U14052 ( .B1(n15079), .B2(n12223), .A(n12222), .ZN(n12224) );
  OAI211_X1 U14053 ( .C1(n10450), .C2(n12226), .A(n12225), .B(n12224), .ZN(
        n12228) );
  NAND2_X1 U14054 ( .A1(n12228), .A2(n15102), .ZN(n12227) );
  OAI21_X1 U14055 ( .B1(n15102), .B2(n8779), .A(n12227), .ZN(P2_U3463) );
  NAND2_X1 U14056 ( .A1(n12228), .A2(n7433), .ZN(n12229) );
  OAI21_X1 U14057 ( .B1(n7433), .B2(n10373), .A(n12229), .ZN(P2_U3510) );
  OAI21_X1 U14058 ( .B1(n12231), .B2(n16556), .A(n12230), .ZN(n12233) );
  AOI211_X1 U14059 ( .C1(n16564), .C2(n12234), .A(n12233), .B(n12232), .ZN(
        n12237) );
  INV_X1 U14060 ( .A(n16469), .ZN(n16565) );
  NAND2_X1 U14061 ( .A1(n16565), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n12235) );
  OAI21_X1 U14062 ( .B1(n12237), .B2(n16565), .A(n12235), .ZN(P1_U3540) );
  NAND2_X1 U14063 ( .A1(n16567), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n12236) );
  OAI21_X1 U14064 ( .B1(n12237), .B2(n16567), .A(n12236), .ZN(P1_U3495) );
  OR2_X1 U14065 ( .A1(n12238), .A2(n12932), .ZN(n12239) );
  NAND2_X1 U14066 ( .A1(n7607), .A2(n12239), .ZN(n12254) );
  OAI22_X1 U14067 ( .A1(n12388), .A2(n13970), .B1(n12544), .B2(n13880), .ZN(
        n12245) );
  NAND2_X1 U14068 ( .A1(n12241), .A2(n12932), .ZN(n12242) );
  AOI21_X1 U14069 ( .B1(n12243), .B2(n12242), .A(n13878), .ZN(n12244) );
  AOI211_X1 U14070 ( .C1(n14052), .C2(n12254), .A(n12245), .B(n12244), .ZN(
        n12256) );
  AOI22_X1 U14071 ( .A1(n13910), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n13980), 
        .B2(n12392), .ZN(n12246) );
  OAI21_X1 U14072 ( .B1(n12823), .B2(n13940), .A(n12246), .ZN(n12247) );
  AOI21_X1 U14073 ( .B1(n12254), .B2(n13846), .A(n12247), .ZN(n12248) );
  OAI21_X1 U14074 ( .B1(n12256), .B2(n13958), .A(n12248), .ZN(P3_U3225) );
  OAI22_X1 U14075 ( .A1(n14051), .A2(n12823), .B1(n16587), .B2(n12249), .ZN(
        n12250) );
  AOI21_X1 U14076 ( .B1(n12254), .B2(n16539), .A(n12250), .ZN(n12251) );
  OAI21_X1 U14077 ( .B1(n12256), .B2(n16585), .A(n12251), .ZN(P3_U3467) );
  INV_X1 U14078 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n12252) );
  OAI22_X1 U14079 ( .A1(n14139), .A2(n12823), .B1(n16590), .B2(n12252), .ZN(
        n12253) );
  AOI21_X1 U14080 ( .B1(n12254), .B2(n14134), .A(n12253), .ZN(n12255) );
  OAI21_X1 U14081 ( .B1(n12256), .B2(n16588), .A(n12255), .ZN(P3_U3414) );
  INV_X1 U14082 ( .A(n12257), .ZN(n12259) );
  INV_X1 U14083 ( .A(SI_24_), .ZN(n12258) );
  OAI222_X1 U14084 ( .A1(P3_U3151), .A2(n12260), .B1(n14154), .B2(n12259), 
        .C1(n12258), .C2(n14150), .ZN(P3_U3271) );
  AND2_X1 U14085 ( .A1(n16606), .A2(n14724), .ZN(n12261) );
  OR2_X1 U14086 ( .A1(n12263), .A2(n12267), .ZN(n12375) );
  NAND2_X1 U14087 ( .A1(n12263), .A2(n12267), .ZN(n12264) );
  OAI22_X1 U14088 ( .A1(n12571), .A2(n14953), .B1(n12265), .B2(n14951), .ZN(
        n12272) );
  INV_X1 U14089 ( .A(n12267), .ZN(n12269) );
  NAND3_X1 U14090 ( .A1(n12266), .A2(n12269), .A3(n12268), .ZN(n12270) );
  AOI21_X1 U14091 ( .B1(n12371), .B2(n12270), .A(n14949), .ZN(n12271) );
  AOI211_X1 U14092 ( .C1(n16507), .C2(n12425), .A(n12272), .B(n12271), .ZN(
        n12429) );
  AOI211_X1 U14093 ( .C1(n12427), .C2(n12273), .A(n14986), .B(n7560), .ZN(
        n12426) );
  NAND2_X1 U14094 ( .A1(n12426), .A2(n16508), .ZN(n12277) );
  INV_X1 U14095 ( .A(n12274), .ZN(n12275) );
  AOI22_X1 U14096 ( .A1(n14992), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12275), 
        .B2(n16511), .ZN(n12276) );
  OAI211_X1 U14097 ( .C1(n7955), .C2(n16515), .A(n12277), .B(n12276), .ZN(
        n12278) );
  AOI21_X1 U14098 ( .B1(n12425), .B2(n16519), .A(n12278), .ZN(n12279) );
  OAI21_X1 U14099 ( .B1(n12429), .B2(n14992), .A(n12279), .ZN(P2_U3252) );
  MUX2_X1 U14100 ( .A(n12280), .B(n12284), .S(n16587), .Z(n12282) );
  AOI22_X1 U14101 ( .A1(n12283), .A2(n16539), .B1(n13445), .B2(n10089), .ZN(
        n12281) );
  NAND2_X1 U14102 ( .A1(n12282), .A2(n12281), .ZN(P3_U3466) );
  INV_X1 U14103 ( .A(n12283), .ZN(n12288) );
  MUX2_X1 U14104 ( .A(n12285), .B(n12284), .S(n13977), .Z(n12287) );
  AOI22_X1 U14105 ( .A1(n13981), .A2(n13445), .B1(n13980), .B2(n13446), .ZN(
        n12286) );
  OAI211_X1 U14106 ( .C1(n12288), .C2(n13984), .A(n12287), .B(n12286), .ZN(
        P3_U3226) );
  INV_X1 U14107 ( .A(n12829), .ZN(n12289) );
  XNOR2_X1 U14108 ( .A(n12290), .B(n7461), .ZN(n16538) );
  XNOR2_X1 U14109 ( .A(n12291), .B(n7461), .ZN(n12293) );
  AOI22_X1 U14110 ( .A1(n13954), .A2(n13604), .B1(n12832), .B2(n13967), .ZN(
        n12292) );
  OAI21_X1 U14111 ( .B1(n12293), .B2(n13878), .A(n12292), .ZN(n12294) );
  AOI21_X1 U14112 ( .B1(n16538), .B2(n14052), .A(n12294), .ZN(n12422) );
  AOI22_X1 U14113 ( .A1(n13910), .A2(P3_REG2_REG_9__SCAN_IN), .B1(n13980), 
        .B2(n12453), .ZN(n12295) );
  OAI21_X1 U14114 ( .B1(n12462), .B2(n13940), .A(n12295), .ZN(n12296) );
  AOI21_X1 U14115 ( .B1(n16538), .B2(n13846), .A(n12296), .ZN(n12297) );
  OAI21_X1 U14116 ( .B1(n12422), .B2(n13958), .A(n12297), .ZN(P3_U3224) );
  OAI222_X1 U14117 ( .A1(n15131), .A2(n12299), .B1(n9157), .B2(P2_U3088), .C1(
        n12298), .C2(n15133), .ZN(P2_U3305) );
  AOI21_X1 U14118 ( .B1(n12300), .B2(n12934), .A(n13878), .ZN(n12303) );
  OAI22_X1 U14119 ( .A1(n13971), .A2(n13880), .B1(n12544), .B2(n13970), .ZN(
        n12301) );
  AOI21_X1 U14120 ( .B1(n12303), .B2(n12302), .A(n12301), .ZN(n12529) );
  INV_X1 U14121 ( .A(n12304), .ZN(n12556) );
  OAI22_X1 U14122 ( .A1(n13977), .A2(n11718), .B1(n12556), .B2(n13946), .ZN(
        n12305) );
  AOI21_X1 U14123 ( .B1(n12546), .B2(n13981), .A(n12305), .ZN(n12309) );
  XNOR2_X1 U14124 ( .A(n12307), .B(n12306), .ZN(n12527) );
  NAND2_X1 U14125 ( .A1(n12527), .A2(n13942), .ZN(n12308) );
  OAI211_X1 U14126 ( .C1(n12529), .C2(n13910), .A(n12309), .B(n12308), .ZN(
        P3_U3223) );
  OR2_X1 U14127 ( .A1(n15940), .A2(n12359), .ZN(n12310) );
  NAND2_X1 U14128 ( .A1(n12312), .A2(n13289), .ZN(n12315) );
  AOI22_X1 U14129 ( .A1(n13155), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n12313), 
        .B2(n13154), .ZN(n12314) );
  XNOR2_X1 U14130 ( .A(n13102), .B(n15371), .ZN(n13329) );
  XNOR2_X1 U14131 ( .A(n12409), .B(n13329), .ZN(n15937) );
  OR2_X1 U14132 ( .A1(n15940), .A2(n15372), .ZN(n12316) );
  INV_X1 U14133 ( .A(n12407), .ZN(n12318) );
  AOI21_X1 U14134 ( .B1(n13329), .B2(n12319), .A(n12318), .ZN(n15935) );
  INV_X1 U14135 ( .A(n13102), .ZN(n15933) );
  NAND2_X1 U14136 ( .A1(n12320), .A2(n15933), .ZN(n12410) );
  OAI211_X1 U14137 ( .C1(n12320), .C2(n15933), .A(n15910), .B(n12410), .ZN(
        n15932) );
  NAND2_X1 U14138 ( .A1(n12321), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n12413) );
  OR2_X1 U14139 ( .A1(n12321), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n12322) );
  NAND2_X1 U14140 ( .A1(n12413), .A2(n12322), .ZN(n15361) );
  NAND2_X1 U14141 ( .A1(n13170), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n12324) );
  NAND2_X1 U14142 ( .A1(n13277), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n12323) );
  AND2_X1 U14143 ( .A1(n12324), .A2(n12323), .ZN(n12327) );
  OR2_X1 U14144 ( .A1(n13284), .A2(n12325), .ZN(n12326) );
  OAI211_X1 U14145 ( .C1(n15361), .C2(n13282), .A(n12327), .B(n12326), .ZN(
        n15540) );
  AOI22_X1 U14146 ( .A1(n15540), .A2(n15789), .B1(n15787), .B2(n15372), .ZN(
        n15931) );
  OAI22_X1 U14147 ( .A1(n16605), .A2(n15931), .B1(n12521), .B2(n16395), .ZN(
        n12329) );
  NOR2_X1 U14148 ( .A1(n15933), .A2(n16595), .ZN(n12328) );
  AOI211_X1 U14149 ( .C1(n16605), .C2(P1_REG2_REG_14__SCAN_IN), .A(n12329), 
        .B(n12328), .ZN(n12330) );
  OAI21_X1 U14150 ( .B1(n15780), .B2(n15932), .A(n12330), .ZN(n12331) );
  AOI21_X1 U14151 ( .B1(n15935), .B2(n15818), .A(n12331), .ZN(n12332) );
  OAI21_X1 U14152 ( .B1(n15821), .B2(n15937), .A(n12332), .ZN(P1_U3279) );
  NAND2_X1 U14153 ( .A1(n12336), .A2(n12335), .ZN(n12338) );
  XNOR2_X1 U14154 ( .A(n13128), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n12337) );
  NAND2_X1 U14155 ( .A1(n12337), .A2(n12338), .ZN(n12576) );
  OAI211_X1 U14156 ( .C1(n12338), .C2(n12337), .A(n15516), .B(n12576), .ZN(
        n12347) );
  NAND2_X1 U14157 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n15297)
         );
  XNOR2_X1 U14158 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n13128), .ZN(n12343) );
  INV_X1 U14159 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n12341) );
  OAI21_X1 U14160 ( .B1(n12341), .B2(n12340), .A(n12339), .ZN(n12342) );
  NAND2_X1 U14161 ( .A1(n12343), .A2(n12342), .ZN(n12579) );
  OAI211_X1 U14162 ( .C1(n12343), .C2(n12342), .A(n15517), .B(n12579), .ZN(
        n12344) );
  NAND2_X1 U14163 ( .A1(n15297), .A2(n12344), .ZN(n12345) );
  AOI21_X1 U14164 ( .B1(n16162), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n12345), 
        .ZN(n12346) );
  OAI211_X1 U14165 ( .C1(n15511), .C2(n13128), .A(n12347), .B(n12346), .ZN(
        P1_U3260) );
  OAI222_X1 U14166 ( .A1(n14154), .A2(n12350), .B1(n14150), .B2(n12349), .C1(
        P3_U3151), .C2(n12348), .ZN(P3_U3270) );
  INV_X1 U14167 ( .A(n12351), .ZN(n12353) );
  OR2_X1 U14168 ( .A1(n12353), .A2(n12352), .ZN(n12354) );
  NAND2_X1 U14169 ( .A1(n12355), .A2(n12354), .ZN(n12362) );
  NAND2_X1 U14170 ( .A1(n15940), .A2(n15255), .ZN(n12357) );
  NAND2_X1 U14171 ( .A1(n15372), .A2(n7432), .ZN(n12356) );
  NAND2_X1 U14172 ( .A1(n12357), .A2(n12356), .ZN(n12358) );
  XNOR2_X1 U14173 ( .A(n12358), .B(n15253), .ZN(n12514) );
  NOR2_X1 U14174 ( .A1(n12359), .A2(n15223), .ZN(n12360) );
  AOI21_X1 U14175 ( .B1(n15940), .B2(n7432), .A(n12360), .ZN(n12512) );
  XNOR2_X1 U14176 ( .A(n12514), .B(n12512), .ZN(n12361) );
  OAI211_X1 U14177 ( .C1(n12362), .C2(n12361), .A(n12516), .B(n15332), .ZN(
        n12367) );
  OAI22_X1 U14178 ( .A1(n15362), .A2(n15358), .B1(n12363), .B2(n15360), .ZN(
        n12364) );
  AOI211_X1 U14179 ( .C1(n15337), .C2(n15373), .A(n12365), .B(n12364), .ZN(
        n12366) );
  OAI211_X1 U14180 ( .C1(n12368), .C2(n15340), .A(n12367), .B(n12366), .ZN(
        P1_U3234) );
  NAND2_X1 U14181 ( .A1(n12427), .A2(n12369), .ZN(n12370) );
  NAND2_X1 U14182 ( .A1(n12371), .A2(n12370), .ZN(n12565) );
  XNOR2_X1 U14183 ( .A(n12565), .B(n12376), .ZN(n12373) );
  OAI21_X1 U14184 ( .B1(n12373), .B2(n14949), .A(n12372), .ZN(n16618) );
  INV_X1 U14185 ( .A(n16618), .ZN(n12383) );
  NAND2_X1 U14186 ( .A1(n12427), .A2(n14723), .ZN(n12374) );
  OAI21_X1 U14187 ( .B1(n12377), .B2(n12376), .A(n12558), .ZN(n16620) );
  OAI211_X1 U14188 ( .C1(n7560), .C2(n16617), .A(n14930), .B(n12560), .ZN(
        n16615) );
  AOI22_X1 U14189 ( .A1(n14992), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n12378), 
        .B2(n16511), .ZN(n12380) );
  NAND2_X1 U14190 ( .A1(n12566), .A2(n16419), .ZN(n12379) );
  OAI211_X1 U14191 ( .C1(n16615), .C2(n14926), .A(n12380), .B(n12379), .ZN(
        n12381) );
  AOI21_X1 U14192 ( .B1(n16620), .B2(n16417), .A(n12381), .ZN(n12382) );
  OAI21_X1 U14193 ( .B1(n12383), .B2(n14992), .A(n12382), .ZN(P2_U3251) );
  XNOR2_X1 U14194 ( .A(n12395), .B(n13428), .ZN(n12454) );
  XNOR2_X1 U14195 ( .A(n12454), .B(n13604), .ZN(n12456) );
  NAND2_X1 U14196 ( .A1(n12387), .A2(n12386), .ZN(n13440) );
  XNOR2_X1 U14197 ( .A(n13445), .B(n13428), .ZN(n12389) );
  XNOR2_X1 U14198 ( .A(n12389), .B(n12394), .ZN(n13441) );
  NAND2_X1 U14199 ( .A1(n13440), .A2(n13441), .ZN(n12391) );
  NAND2_X1 U14200 ( .A1(n12391), .A2(n12390), .ZN(n12457) );
  XOR2_X1 U14201 ( .A(n12456), .B(n12457), .Z(n12400) );
  INV_X1 U14202 ( .A(n12392), .ZN(n12398) );
  AOI21_X1 U14203 ( .B1(n12394), .B2(n13589), .A(n12393), .ZN(n12397) );
  AOI22_X1 U14204 ( .A1(n13603), .A2(n13566), .B1(n13596), .B2(n12395), .ZN(
        n12396) );
  OAI211_X1 U14205 ( .C1(n12398), .C2(n13448), .A(n12397), .B(n12396), .ZN(
        n12399) );
  AOI21_X1 U14206 ( .B1(n12400), .B2(n13576), .A(n12399), .ZN(n12401) );
  INV_X1 U14207 ( .A(n12401), .ZN(P3_U3161) );
  NAND2_X1 U14208 ( .A1(n12402), .A2(n13289), .ZN(n12405) );
  AOI22_X1 U14209 ( .A1(n13154), .A2(n12403), .B1(n13155), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n12404) );
  XNOR2_X1 U14210 ( .A(n15561), .B(n15540), .ZN(n15559) );
  NAND2_X1 U14211 ( .A1(n13102), .A2(n15371), .ZN(n12406) );
  XOR2_X1 U14212 ( .A(n15559), .B(n15541), .Z(n15930) );
  NAND2_X1 U14213 ( .A1(n13102), .A2(n15358), .ZN(n12408) );
  XOR2_X1 U14214 ( .A(n15559), .B(n15560), .Z(n15928) );
  AOI21_X1 U14215 ( .B1(n12410), .B2(n15561), .A(n15915), .ZN(n12411) );
  NAND2_X1 U14216 ( .A1(n12411), .A2(n15802), .ZN(n15925) );
  INV_X1 U14217 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n12412) );
  NAND2_X1 U14218 ( .A1(n12413), .A2(n12412), .ZN(n12414) );
  NAND2_X1 U14219 ( .A1(n13122), .A2(n12414), .ZN(n15804) );
  AOI22_X1 U14220 ( .A1(n13170), .A2(P1_REG0_REG_16__SCAN_IN), .B1(n13277), 
        .B2(P1_REG2_REG_16__SCAN_IN), .ZN(n12416) );
  NAND2_X1 U14221 ( .A1(n8317), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n12415) );
  OAI211_X1 U14222 ( .C1(n15804), .C2(n13282), .A(n12416), .B(n12415), .ZN(
        n15788) );
  AOI22_X1 U14223 ( .A1(n15788), .A2(n15789), .B1(n15787), .B2(n15371), .ZN(
        n15924) );
  OAI22_X1 U14224 ( .A1(n16605), .A2(n15924), .B1(n15361), .B2(n16395), .ZN(
        n12418) );
  INV_X1 U14225 ( .A(n15561), .ZN(n15926) );
  NOR2_X1 U14226 ( .A1(n15926), .A2(n16595), .ZN(n12417) );
  AOI211_X1 U14227 ( .C1(n16605), .C2(P1_REG2_REG_15__SCAN_IN), .A(n12418), 
        .B(n12417), .ZN(n12419) );
  OAI21_X1 U14228 ( .B1(n15780), .B2(n15925), .A(n12419), .ZN(n12420) );
  AOI21_X1 U14229 ( .B1(n15928), .B2(n15711), .A(n12420), .ZN(n12421) );
  OAI21_X1 U14230 ( .B1(n15930), .B2(n16597), .A(n12421), .ZN(P1_U3278) );
  OAI21_X1 U14231 ( .B1(n12462), .B2(n16580), .A(n12422), .ZN(n16540) );
  INV_X1 U14232 ( .A(n16540), .ZN(n12424) );
  AOI22_X1 U14233 ( .A1(n16538), .A2(n14134), .B1(P3_REG0_REG_9__SCAN_IN), 
        .B2(n16588), .ZN(n12423) );
  OAI21_X1 U14234 ( .B1(n12424), .B2(n16588), .A(n12423), .ZN(P3_U3417) );
  INV_X1 U14235 ( .A(n12425), .ZN(n12430) );
  AOI21_X1 U14236 ( .B1(n15079), .B2(n12427), .A(n12426), .ZN(n12428) );
  OAI211_X1 U14237 ( .C1(n10450), .C2(n12430), .A(n12429), .B(n12428), .ZN(
        n12433) );
  NAND2_X1 U14238 ( .A1(n12433), .A2(n7433), .ZN(n12431) );
  OAI21_X1 U14239 ( .B1(n7433), .B2(n12432), .A(n12431), .ZN(P2_U3512) );
  NAND2_X1 U14240 ( .A1(n12433), .A2(n15102), .ZN(n12434) );
  OAI21_X1 U14241 ( .B1(n15102), .B2(n8817), .A(n12434), .ZN(P2_U3469) );
  INV_X1 U14242 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12437) );
  AOI21_X1 U14243 ( .B1(n12437), .B2(n12436), .A(n12487), .ZN(n12452) );
  XNOR2_X1 U14244 ( .A(n12492), .B(n12486), .ZN(n12439) );
  NAND2_X1 U14245 ( .A1(P3_REG2_REG_13__SCAN_IN), .A2(n12439), .ZN(n12493) );
  OAI21_X1 U14246 ( .B1(P3_REG2_REG_13__SCAN_IN), .B2(n12439), .A(n12493), 
        .ZN(n12450) );
  NOR2_X1 U14247 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14493), .ZN(n13548) );
  AOI21_X1 U14248 ( .B1(n16036), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n13548), 
        .ZN(n12440) );
  OAI21_X1 U14249 ( .B1(n16367), .B2(n12498), .A(n12440), .ZN(n12449) );
  MUX2_X1 U14250 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n7429), .Z(n12499) );
  XNOR2_X1 U14251 ( .A(n12499), .B(n12498), .ZN(n12446) );
  MUX2_X1 U14252 ( .A(n12442), .B(n12441), .S(n7429), .Z(n12443) );
  NAND2_X1 U14253 ( .A1(n12444), .A2(n12443), .ZN(n12445) );
  NOR2_X1 U14254 ( .A1(n12445), .A2(n12446), .ZN(n12501) );
  AOI21_X1 U14255 ( .B1(n12446), .B2(n12445), .A(n12501), .ZN(n12447) );
  NOR2_X1 U14256 ( .A1(n12447), .A2(n16376), .ZN(n12448) );
  AOI211_X1 U14257 ( .C1(n13712), .C2(n12450), .A(n12449), .B(n12448), .ZN(
        n12451) );
  OAI21_X1 U14258 ( .B1(n12452), .B2(n16374), .A(n12451), .ZN(P3_U3195) );
  INV_X1 U14259 ( .A(n12453), .ZN(n12467) );
  XNOR2_X1 U14260 ( .A(n12462), .B(n13428), .ZN(n12543) );
  XNOR2_X1 U14261 ( .A(n12543), .B(n12544), .ZN(n12459) );
  INV_X1 U14262 ( .A(n12454), .ZN(n12455) );
  OAI21_X1 U14263 ( .B1(n12459), .B2(n12458), .A(n12549), .ZN(n12460) );
  NAND2_X1 U14264 ( .A1(n12460), .A2(n13576), .ZN(n12466) );
  OAI22_X1 U14265 ( .A1(n13582), .A2(n12462), .B1(n12461), .B2(n13593), .ZN(
        n12463) );
  AOI211_X1 U14266 ( .C1(n13589), .C2(n13604), .A(n12464), .B(n12463), .ZN(
        n12465) );
  OAI211_X1 U14267 ( .C1(n12467), .C2(n13448), .A(n12466), .B(n12465), .ZN(
        P3_U3171) );
  INV_X1 U14268 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n13219) );
  NAND2_X1 U14269 ( .A1(n13218), .A2(n12468), .ZN(n12469) );
  OAI211_X1 U14270 ( .C1(n13219), .C2(n15987), .A(n12469), .B(n13369), .ZN(
        P1_U3332) );
  NAND2_X1 U14271 ( .A1(n13218), .A2(n12470), .ZN(n12472) );
  OAI211_X1 U14272 ( .C1(n12473), .C2(n15133), .A(n12472), .B(n12471), .ZN(
        P2_U3304) );
  XNOR2_X1 U14273 ( .A(n12474), .B(n12936), .ZN(n16579) );
  INV_X1 U14274 ( .A(n16579), .ZN(n12482) );
  XNOR2_X1 U14275 ( .A(n12475), .B(n12936), .ZN(n12476) );
  NAND2_X1 U14276 ( .A1(n12476), .A2(n13973), .ZN(n12478) );
  AOI22_X1 U14277 ( .A1(n13954), .A2(n12832), .B1(n13953), .B2(n13967), .ZN(
        n12477) );
  NAND2_X1 U14278 ( .A1(n12478), .A2(n12477), .ZN(n16582) );
  AOI22_X1 U14279 ( .A1(n13910), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n13980), 
        .B2(n12661), .ZN(n12479) );
  OAI21_X1 U14280 ( .B1(n16581), .B2(n13940), .A(n12479), .ZN(n12480) );
  AOI21_X1 U14281 ( .B1(n16582), .B2(n13977), .A(n12480), .ZN(n12481) );
  OAI21_X1 U14282 ( .B1(n13963), .B2(n12482), .A(n12481), .ZN(P3_U3222) );
  INV_X1 U14283 ( .A(SI_26_), .ZN(n12484) );
  OAI222_X1 U14284 ( .A1(n14154), .A2(n8177), .B1(n14150), .B2(n12484), .C1(
        P3_U3151), .C2(n12483), .ZN(P3_U3269) );
  NAND2_X1 U14285 ( .A1(n13618), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13608) );
  INV_X1 U14286 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n14049) );
  NAND2_X1 U14287 ( .A1(n13628), .A2(n14049), .ZN(n12488) );
  NAND2_X1 U14288 ( .A1(n13608), .A2(n12488), .ZN(n12490) );
  INV_X1 U14289 ( .A(n13609), .ZN(n12489) );
  AOI21_X1 U14290 ( .B1(n12491), .B2(n12490), .A(n12489), .ZN(n12507) );
  NAND2_X1 U14291 ( .A1(n12498), .A2(n12492), .ZN(n12494) );
  XNOR2_X1 U14292 ( .A(P3_REG2_REG_14__SCAN_IN), .B(n13618), .ZN(n12495) );
  XNOR2_X1 U14293 ( .A(n13631), .B(n12495), .ZN(n12497) );
  NOR2_X1 U14294 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n14464), .ZN(n13464) );
  AOI21_X1 U14295 ( .B1(n16036), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n13464), 
        .ZN(n12496) );
  OAI21_X1 U14296 ( .B1(n16382), .B2(n12497), .A(n12496), .ZN(n12505) );
  MUX2_X1 U14297 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n7429), .Z(n13619) );
  XOR2_X1 U14298 ( .A(n13628), .B(n13619), .Z(n12503) );
  NOR2_X1 U14299 ( .A1(n12499), .A2(n12498), .ZN(n12500) );
  OR2_X1 U14300 ( .A1(n12501), .A2(n12500), .ZN(n12502) );
  AOI211_X1 U14301 ( .C1(n12503), .C2(n12502), .A(n16376), .B(n13617), .ZN(
        n12504) );
  AOI211_X1 U14302 ( .C1(n13707), .C2(n13628), .A(n12505), .B(n12504), .ZN(
        n12506) );
  OAI21_X1 U14303 ( .B1(n12507), .B2(n16374), .A(n12506), .ZN(P3_U3196) );
  NAND2_X1 U14304 ( .A1(n13102), .A2(n15255), .ZN(n12509) );
  NAND2_X1 U14305 ( .A1(n15371), .A2(n7432), .ZN(n12508) );
  NAND2_X1 U14306 ( .A1(n12509), .A2(n12508), .ZN(n12510) );
  XNOR2_X1 U14307 ( .A(n12510), .B(n15221), .ZN(n15146) );
  AND2_X1 U14308 ( .A1(n15252), .A2(n15371), .ZN(n12511) );
  AOI21_X1 U14309 ( .B1(n13102), .B2(n7432), .A(n12511), .ZN(n15145) );
  XNOR2_X1 U14310 ( .A(n15146), .B(n15145), .ZN(n12520) );
  INV_X1 U14311 ( .A(n12512), .ZN(n12513) );
  NAND2_X1 U14312 ( .A1(n12514), .A2(n12513), .ZN(n12515) );
  INV_X1 U14313 ( .A(n15148), .ZN(n12518) );
  AOI21_X1 U14314 ( .B1(n12520), .B2(n12519), .A(n12518), .ZN(n12526) );
  NOR2_X1 U14315 ( .A1(n15360), .A2(n12521), .ZN(n12524) );
  OAI21_X1 U14316 ( .B1(n15931), .B2(n15264), .A(n12522), .ZN(n12523) );
  AOI211_X1 U14317 ( .C1(n13102), .C2(n15365), .A(n12524), .B(n12523), .ZN(
        n12525) );
  OAI21_X1 U14318 ( .B1(n12526), .B2(n15367), .A(n12525), .ZN(P1_U3215) );
  INV_X1 U14319 ( .A(n12546), .ZN(n12833) );
  INV_X1 U14320 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n12530) );
  NAND2_X1 U14321 ( .A1(n12527), .A2(n16578), .ZN(n12528) );
  AND2_X1 U14322 ( .A1(n12529), .A2(n12528), .ZN(n12532) );
  MUX2_X1 U14323 ( .A(n12530), .B(n12532), .S(n16590), .Z(n12531) );
  OAI21_X1 U14324 ( .B1(n14139), .B2(n12833), .A(n12531), .ZN(P3_U3420) );
  MUX2_X1 U14325 ( .A(n11733), .B(n12532), .S(n16587), .Z(n12533) );
  OAI21_X1 U14326 ( .B1(n14051), .B2(n12833), .A(n12533), .ZN(P3_U3469) );
  NOR2_X1 U14327 ( .A1(n14683), .A2(n12654), .ZN(n12536) );
  AOI22_X1 U14328 ( .A1(n14718), .A2(n14913), .B1(n14911), .B2(n14720), .ZN(
        n12646) );
  OAI22_X1 U14329 ( .A1(n14650), .A2(n12646), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12534), .ZN(n12535) );
  AOI211_X1 U14330 ( .C1(n15068), .C2(n14691), .A(n12536), .B(n12535), .ZN(
        n12541) );
  INV_X1 U14331 ( .A(n14720), .ZN(n12640) );
  OAI22_X1 U14332 ( .A1(n12538), .A2(n14686), .B1(n12640), .B2(n14694), .ZN(
        n12539) );
  NAND3_X1 U14333 ( .A1(n12634), .A2(n8040), .A3(n12539), .ZN(n12540) );
  OAI211_X1 U14334 ( .C1(n12542), .C2(n14686), .A(n12541), .B(n12540), .ZN(
        P2_U3200) );
  INV_X1 U14335 ( .A(n12543), .ZN(n12545) );
  NAND2_X1 U14336 ( .A1(n12545), .A2(n12544), .ZN(n12547) );
  AND2_X1 U14337 ( .A1(n12549), .A2(n12547), .ZN(n12551) );
  XNOR2_X1 U14338 ( .A(n12546), .B(n13428), .ZN(n12613) );
  XNOR2_X1 U14339 ( .A(n12613), .B(n12832), .ZN(n12550) );
  OAI211_X1 U14340 ( .C1(n12551), .C2(n12550), .A(n13576), .B(n12616), .ZN(
        n12555) );
  OAI22_X1 U14341 ( .A1(n13582), .A2(n12833), .B1(n13971), .B2(n13593), .ZN(
        n12552) );
  AOI211_X1 U14342 ( .C1(n13589), .C2(n13603), .A(n12553), .B(n12552), .ZN(
        n12554) );
  OAI211_X1 U14343 ( .C1(n12556), .C2(n13448), .A(n12555), .B(n12554), .ZN(
        P3_U3157) );
  OR2_X1 U14344 ( .A1(n12566), .A2(n14722), .ZN(n12557) );
  NAND2_X1 U14345 ( .A1(n12558), .A2(n12557), .ZN(n12591) );
  XNOR2_X1 U14346 ( .A(n12591), .B(n12569), .ZN(n15083) );
  OR2_X1 U14347 ( .A1(n12560), .A2(n15078), .ZN(n12595) );
  INV_X1 U14348 ( .A(n12595), .ZN(n12559) );
  AOI211_X1 U14349 ( .C1(n15078), .C2(n12560), .A(n14986), .B(n12559), .ZN(
        n15077) );
  INV_X1 U14350 ( .A(n15078), .ZN(n12563) );
  INV_X1 U14351 ( .A(n12606), .ZN(n12561) );
  AOI22_X1 U14352 ( .A1(n16522), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n12561), 
        .B2(n16511), .ZN(n12562) );
  OAI21_X1 U14353 ( .B1(n12563), .B2(n16515), .A(n12562), .ZN(n12574) );
  OR2_X1 U14354 ( .A1(n12566), .A2(n12571), .ZN(n12564) );
  NAND2_X1 U14355 ( .A1(n12565), .A2(n12564), .ZN(n12568) );
  NAND2_X1 U14356 ( .A1(n12566), .A2(n12571), .ZN(n12567) );
  INV_X1 U14357 ( .A(n12569), .ZN(n12590) );
  AOI21_X1 U14358 ( .B1(n12570), .B2(n12590), .A(n14949), .ZN(n12572) );
  OAI22_X1 U14359 ( .A1(n12640), .A2(n14953), .B1(n12571), .B2(n14951), .ZN(
        n12604) );
  AOI21_X1 U14360 ( .B1(n12572), .B2(n12587), .A(n12604), .ZN(n15081) );
  NOR2_X1 U14361 ( .A1(n15081), .A2(n14992), .ZN(n12573) );
  AOI211_X1 U14362 ( .C1(n15077), .C2(n16508), .A(n12574), .B(n12573), .ZN(
        n12575) );
  OAI21_X1 U14363 ( .B1(n14892), .B2(n15083), .A(n12575), .ZN(P2_U3250) );
  INV_X1 U14364 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n12577) );
  OAI21_X1 U14365 ( .B1(n12577), .B2(n13128), .A(n12576), .ZN(n15506) );
  XNOR2_X1 U14366 ( .A(n12585), .B(n15506), .ZN(n12578) );
  NAND2_X1 U14367 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n12578), .ZN(n15508) );
  OAI211_X1 U14368 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n12578), .A(n15516), 
        .B(n15508), .ZN(n12584) );
  NAND2_X1 U14369 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15334)
         );
  INV_X1 U14370 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n13124) );
  XNOR2_X1 U14371 ( .A(n15501), .B(n12585), .ZN(n12580) );
  NAND2_X1 U14372 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n12580), .ZN(n15502) );
  OAI211_X1 U14373 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n12580), .A(n15517), 
        .B(n15502), .ZN(n12581) );
  NAND2_X1 U14374 ( .A1(n15334), .A2(n12581), .ZN(n12582) );
  AOI21_X1 U14375 ( .B1(n16162), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n12582), 
        .ZN(n12583) );
  OAI211_X1 U14376 ( .C1(n15511), .C2(n12585), .A(n12584), .B(n12583), .ZN(
        P1_U3261) );
  OR2_X1 U14377 ( .A1(n15078), .A2(n12626), .ZN(n12586) );
  OAI211_X1 U14378 ( .C1(n12594), .C2(n12588), .A(n12644), .B(n14981), .ZN(
        n12589) );
  AOI22_X1 U14379 ( .A1(n14719), .A2(n14913), .B1(n14911), .B2(n14721), .ZN(
        n12630) );
  AND2_X1 U14380 ( .A1(n12589), .A2(n12630), .ZN(n15075) );
  NAND2_X1 U14381 ( .A1(n12591), .A2(n12590), .ZN(n12593) );
  OR2_X1 U14382 ( .A1(n15078), .A2(n14721), .ZN(n12592) );
  OAI21_X1 U14383 ( .B1(n7547), .B2(n8118), .A(n12649), .ZN(n15076) );
  INV_X1 U14384 ( .A(n15076), .ZN(n12602) );
  INV_X1 U14385 ( .A(n15073), .ZN(n12600) );
  AOI21_X1 U14386 ( .B1(n15073), .B2(n12595), .A(n14986), .ZN(n12596) );
  AND2_X1 U14387 ( .A1(n12651), .A2(n12596), .ZN(n15072) );
  NAND2_X1 U14388 ( .A1(n15072), .A2(n16508), .ZN(n12599) );
  INV_X1 U14389 ( .A(n12633), .ZN(n12597) );
  AOI22_X1 U14390 ( .A1(n14992), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n12597), 
        .B2(n16511), .ZN(n12598) );
  OAI211_X1 U14391 ( .C1(n12600), .C2(n16515), .A(n12599), .B(n12598), .ZN(
        n12601) );
  AOI21_X1 U14392 ( .B1(n12602), .B2(n16417), .A(n12601), .ZN(n12603) );
  OAI21_X1 U14393 ( .B1(n14992), .B2(n15075), .A(n12603), .ZN(P2_U3249) );
  AOI22_X1 U14394 ( .A1(n14681), .A2(n12604), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12605) );
  OAI21_X1 U14395 ( .B1(n12606), .B2(n14683), .A(n12605), .ZN(n12611) );
  INV_X1 U14396 ( .A(n12607), .ZN(n12629) );
  AOI211_X1 U14397 ( .C1(n12609), .C2(n12608), .A(n14686), .B(n12629), .ZN(
        n12610) );
  AOI211_X1 U14398 ( .C1(n15078), .C2(n14691), .A(n12611), .B(n12610), .ZN(
        n12612) );
  INV_X1 U14399 ( .A(n12612), .ZN(P2_U3213) );
  INV_X1 U14400 ( .A(n12613), .ZN(n12614) );
  NAND2_X1 U14401 ( .A1(n12614), .A2(n12832), .ZN(n12615) );
  XNOR2_X1 U14402 ( .A(n16581), .B(n13428), .ZN(n12617) );
  XNOR2_X1 U14403 ( .A(n12617), .B(n13971), .ZN(n12666) );
  XNOR2_X1 U14404 ( .A(n14060), .B(n13428), .ZN(n13377) );
  XNOR2_X1 U14405 ( .A(n13377), .B(n13953), .ZN(n12619) );
  XNOR2_X1 U14406 ( .A(n13374), .B(n12619), .ZN(n12625) );
  NOR2_X1 U14407 ( .A1(n13582), .A2(n14138), .ZN(n12623) );
  NAND2_X1 U14408 ( .A1(n13566), .A2(n13968), .ZN(n12620) );
  OAI211_X1 U14409 ( .C1(n13971), .C2(n13568), .A(n12621), .B(n12620), .ZN(
        n12622) );
  AOI211_X1 U14410 ( .C1(n13979), .C2(n13590), .A(n12623), .B(n12622), .ZN(
        n12624) );
  OAI21_X1 U14411 ( .B1(n12625), .B2(n13599), .A(n12624), .ZN(P3_U3164) );
  NOR3_X1 U14412 ( .A1(n12627), .A2(n12626), .A3(n14694), .ZN(n12628) );
  AOI21_X1 U14413 ( .B1(n12629), .B2(n14707), .A(n12628), .ZN(n12639) );
  INV_X1 U14414 ( .A(n12630), .ZN(n12631) );
  AOI22_X1 U14415 ( .A1(n14681), .A2(n12631), .B1(P2_REG3_REG_16__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12632) );
  OAI21_X1 U14416 ( .B1(n12633), .B2(n14683), .A(n12632), .ZN(n12636) );
  NOR2_X1 U14417 ( .A1(n12634), .A2(n14686), .ZN(n12635) );
  AOI211_X1 U14418 ( .C1(n15073), .C2(n14691), .A(n12636), .B(n12635), .ZN(
        n12637) );
  OAI21_X1 U14419 ( .B1(n12639), .B2(n12638), .A(n12637), .ZN(P2_U3198) );
  OR2_X1 U14420 ( .A1(n15073), .A2(n12640), .ZN(n12643) );
  NAND2_X1 U14421 ( .A1(n12644), .A2(n12643), .ZN(n12641) );
  INV_X1 U14422 ( .A(n12642), .ZN(n12650) );
  NAND3_X1 U14423 ( .A1(n12644), .A2(n12650), .A3(n12643), .ZN(n12645) );
  NAND3_X1 U14424 ( .A1(n12674), .A2(n14981), .A3(n12645), .ZN(n12647) );
  NAND2_X1 U14425 ( .A1(n15073), .A2(n14720), .ZN(n12648) );
  OAI21_X1 U14426 ( .B1(n7557), .B2(n12650), .A(n12698), .ZN(n15066) );
  INV_X1 U14427 ( .A(n15068), .ZN(n12658) );
  NAND2_X1 U14428 ( .A1(n15068), .A2(n12651), .ZN(n12652) );
  NAND2_X1 U14429 ( .A1(n12652), .A2(n14930), .ZN(n12653) );
  NOR2_X1 U14430 ( .A1(n14985), .A2(n12653), .ZN(n15067) );
  NAND2_X1 U14431 ( .A1(n15067), .A2(n16508), .ZN(n12657) );
  INV_X1 U14432 ( .A(n12654), .ZN(n12655) );
  AOI22_X1 U14433 ( .A1(n14992), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n12655), 
        .B2(n16511), .ZN(n12656) );
  OAI211_X1 U14434 ( .C1(n12658), .C2(n16515), .A(n12657), .B(n12656), .ZN(
        n12659) );
  AOI21_X1 U14435 ( .B1(n15066), .B2(n16417), .A(n12659), .ZN(n12660) );
  OAI21_X1 U14436 ( .B1(n14992), .B2(n15070), .A(n12660), .ZN(P2_U3248) );
  INV_X1 U14437 ( .A(n12661), .ZN(n12665) );
  AOI21_X1 U14438 ( .B1(n12832), .B2(n13589), .A(n12662), .ZN(n12664) );
  NAND2_X1 U14439 ( .A1(n13566), .A2(n13953), .ZN(n12663) );
  OAI211_X1 U14440 ( .C1(n13448), .C2(n12665), .A(n12664), .B(n12663), .ZN(
        n12670) );
  XNOR2_X1 U14441 ( .A(n12667), .B(n12666), .ZN(n12668) );
  NOR2_X1 U14442 ( .A1(n12668), .A2(n13599), .ZN(n12669) );
  AOI211_X1 U14443 ( .C1(n13596), .C2(n12671), .A(n12670), .B(n12669), .ZN(
        n12672) );
  INV_X1 U14444 ( .A(n12672), .ZN(P3_U3176) );
  INV_X1 U14445 ( .A(n14719), .ZN(n14680) );
  OR2_X1 U14446 ( .A1(n15068), .A2(n14680), .ZN(n12673) );
  NAND2_X1 U14447 ( .A1(n15062), .A2(n14177), .ZN(n12675) );
  INV_X1 U14448 ( .A(n14717), .ZN(n14950) );
  NOR2_X1 U14449 ( .A1(n15057), .A2(n14950), .ZN(n12677) );
  NAND2_X1 U14450 ( .A1(n15057), .A2(n14950), .ZN(n12676) );
  INV_X1 U14451 ( .A(n14716), .ZN(n14941) );
  AND2_X1 U14452 ( .A1(n15053), .A2(n14941), .ZN(n12678) );
  OR2_X1 U14453 ( .A1(n15053), .A2(n14941), .ZN(n12679) );
  INV_X1 U14454 ( .A(n14912), .ZN(n14952) );
  OR2_X1 U14455 ( .A1(n15048), .A2(n14952), .ZN(n12680) );
  NAND2_X1 U14456 ( .A1(n15039), .A2(n14942), .ZN(n12681) );
  INV_X1 U14457 ( .A(n14914), .ZN(n14648) );
  OR2_X1 U14458 ( .A1(n15035), .A2(n14648), .ZN(n12682) );
  NAND2_X1 U14459 ( .A1(n14896), .A2(n12682), .ZN(n12684) );
  NAND2_X1 U14460 ( .A1(n15035), .A2(n14648), .ZN(n12683) );
  NAND2_X1 U14461 ( .A1(n12684), .A2(n12683), .ZN(n14881) );
  OR2_X1 U14462 ( .A1(n14889), .A2(n14714), .ZN(n12685) );
  NAND2_X1 U14463 ( .A1(n14877), .A2(n14860), .ZN(n12687) );
  NOR2_X1 U14464 ( .A1(n15016), .A2(n14861), .ZN(n14821) );
  NAND2_X1 U14465 ( .A1(n14839), .A2(n14911), .ZN(n12694) );
  INV_X1 U14466 ( .A(P2_B_REG_SCAN_IN), .ZN(n12691) );
  NOR2_X1 U14467 ( .A1(n15119), .A2(n12691), .ZN(n12692) );
  NOR2_X1 U14468 ( .A1(n14953), .A2(n12692), .ZN(n14806) );
  NAND2_X1 U14469 ( .A1(n14806), .A2(n14712), .ZN(n12693) );
  OR2_X1 U14470 ( .A1(n15068), .A2(n14719), .ZN(n12697) );
  NAND2_X1 U14471 ( .A1(n12698), .A2(n12697), .ZN(n14983) );
  NAND2_X1 U14472 ( .A1(n14983), .A2(n14984), .ZN(n12700) );
  NAND2_X1 U14473 ( .A1(n14995), .A2(n14177), .ZN(n12699) );
  NAND2_X1 U14474 ( .A1(n15057), .A2(n14717), .ZN(n12701) );
  OR2_X1 U14475 ( .A1(n14716), .A2(n15053), .ZN(n12702) );
  NAND2_X1 U14476 ( .A1(n14945), .A2(n12702), .ZN(n12704) );
  NAND2_X1 U14477 ( .A1(n15053), .A2(n14716), .ZN(n12703) );
  AND2_X1 U14478 ( .A1(n15048), .A2(n14912), .ZN(n12705) );
  OR2_X2 U14479 ( .A1(n14919), .A2(n7770), .ZN(n15041) );
  NAND2_X1 U14480 ( .A1(n15039), .A2(n14715), .ZN(n12707) );
  OR2_X1 U14481 ( .A1(n15035), .A2(n14914), .ZN(n12708) );
  NAND2_X1 U14482 ( .A1(n15035), .A2(n14914), .ZN(n12709) );
  NAND2_X1 U14483 ( .A1(n14866), .A2(n12710), .ZN(n12712) );
  NAND2_X1 U14484 ( .A1(n12712), .A2(n12711), .ZN(n14851) );
  AND2_X1 U14485 ( .A1(n14856), .A2(n14871), .ZN(n12713) );
  OR2_X1 U14486 ( .A1(n14856), .A2(n14871), .ZN(n12714) );
  INV_X1 U14487 ( .A(n14834), .ZN(n12715) );
  AOI22_X1 U14488 ( .A1(n14818), .A2(n8078), .B1(n14839), .B2(n15011), .ZN(
        n12717) );
  XNOR2_X1 U14489 ( .A(n12717), .B(n12716), .ZN(n15004) );
  INV_X1 U14490 ( .A(n15005), .ZN(n12723) );
  INV_X1 U14491 ( .A(n15039), .ZN(n12719) );
  INV_X1 U14492 ( .A(n15053), .ZN(n14960) );
  NAND2_X1 U14493 ( .A1(n14960), .A2(n12718), .ZN(n14955) );
  NAND2_X1 U14494 ( .A1(n12719), .A2(n14933), .ZN(n14918) );
  OAI211_X1 U14495 ( .C1(n12723), .C2(n14824), .A(n14930), .B(n14811), .ZN(
        n15006) );
  NOR2_X1 U14496 ( .A1(n15006), .A2(n14926), .ZN(n12725) );
  INV_X1 U14497 ( .A(n12720), .ZN(n12721) );
  AOI22_X1 U14498 ( .A1(n12721), .A2(n16511), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14992), .ZN(n12722) );
  OAI21_X1 U14499 ( .B1(n12723), .B2(n16515), .A(n12722), .ZN(n12724) );
  AOI211_X1 U14500 ( .C1(n15004), .C2(n16417), .A(n12725), .B(n12724), .ZN(
        n12726) );
  OAI21_X1 U14501 ( .B1(n15009), .B2(n14992), .A(n12726), .ZN(P2_U3236) );
  OAI222_X1 U14502 ( .A1(n15133), .A2(n12729), .B1(n15123), .B2(n12728), .C1(
        P2_U3088), .C2(n12727), .ZN(P2_U3308) );
  OAI222_X1 U14503 ( .A1(n15131), .A2(n15975), .B1(n12730), .B2(P2_U3088), 
        .C1(n12731), .C2(n15133), .ZN(P2_U3297) );
  OAI222_X1 U14504 ( .A1(n14154), .A2(n12733), .B1(n14150), .B2(n14407), .C1(
        P3_U3151), .C2(n12732), .ZN(P3_U3267) );
  INV_X1 U14505 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12740) );
  NAND2_X1 U14506 ( .A1(n9984), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12738) );
  INV_X1 U14507 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12735) );
  OR2_X1 U14508 ( .A1(n7434), .A2(n12735), .ZN(n12737) );
  OAI211_X1 U14509 ( .C1(n12740), .C2(n7436), .A(n12738), .B(n12737), .ZN(
        n12741) );
  INV_X1 U14510 ( .A(n12741), .ZN(n12742) );
  INV_X1 U14511 ( .A(n12744), .ZN(n12745) );
  NAND2_X1 U14512 ( .A1(n12746), .A2(n12745), .ZN(n12748) );
  NAND2_X1 U14513 ( .A1(n15977), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12747) );
  NAND2_X1 U14514 ( .A1(n12748), .A2(n12747), .ZN(n12754) );
  XNOR2_X1 U14515 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n12753) );
  INV_X1 U14516 ( .A(n12753), .ZN(n12749) );
  XNOR2_X1 U14517 ( .A(n12754), .B(n12749), .ZN(n13436) );
  NAND2_X1 U14518 ( .A1(n13436), .A2(n12759), .ZN(n12751) );
  NAND2_X1 U14519 ( .A1(n12760), .A2(SI_30_), .ZN(n12750) );
  OAI21_X1 U14520 ( .B1(n12913), .B2(n13717), .A(n13720), .ZN(n12752) );
  AND2_X1 U14521 ( .A1(n12752), .A2(n12906), .ZN(n12957) );
  NAND2_X1 U14522 ( .A1(n12754), .A2(n12753), .ZN(n12756) );
  INV_X1 U14523 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n15974) );
  NAND2_X1 U14524 ( .A1(n15974), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12755) );
  NAND2_X1 U14525 ( .A1(n12756), .A2(n12755), .ZN(n12758) );
  XNOR2_X1 U14526 ( .A(n15107), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n12757) );
  XNOR2_X1 U14527 ( .A(n12758), .B(n12757), .ZN(n14142) );
  NAND2_X1 U14528 ( .A1(n14142), .A2(n12759), .ZN(n12762) );
  NAND2_X1 U14529 ( .A1(n12760), .A2(SI_31_), .ZN(n12761) );
  NAND2_X1 U14530 ( .A1(n12762), .A2(n12761), .ZN(n13715) );
  OR2_X1 U14531 ( .A1(n13715), .A2(n13717), .ZN(n12955) );
  OR2_X1 U14532 ( .A1(n13720), .A2(n12913), .ZN(n12914) );
  INV_X1 U14533 ( .A(n13717), .ZN(n13601) );
  NAND2_X1 U14534 ( .A1(n12914), .A2(n13601), .ZN(n12764) );
  NAND2_X1 U14535 ( .A1(n12764), .A2(n13715), .ZN(n12915) );
  XNOR2_X1 U14536 ( .A(n12915), .B(n13694), .ZN(n12765) );
  NAND2_X1 U14537 ( .A1(n12771), .A2(n12769), .ZN(n13764) );
  INV_X1 U14538 ( .A(n13777), .ZN(n12766) );
  NAND2_X1 U14539 ( .A1(n12767), .A2(n13750), .ZN(n12947) );
  INV_X1 U14540 ( .A(n12781), .ZN(n12776) );
  NAND2_X1 U14541 ( .A1(n12769), .A2(n12768), .ZN(n12770) );
  NAND3_X1 U14542 ( .A1(n12772), .A2(n12771), .A3(n12770), .ZN(n12774) );
  NAND2_X1 U14543 ( .A1(n13759), .A2(n13733), .ZN(n12773) );
  NAND2_X1 U14544 ( .A1(n12774), .A2(n12773), .ZN(n12777) );
  INV_X1 U14545 ( .A(n12777), .ZN(n12775) );
  OAI21_X1 U14546 ( .B1(n12947), .B2(n12776), .A(n12775), .ZN(n12779) );
  INV_X1 U14547 ( .A(n12780), .ZN(n12778) );
  INV_X1 U14548 ( .A(n12782), .ZN(n12783) );
  NAND2_X1 U14549 ( .A1(n12784), .A2(n12783), .ZN(n12786) );
  NAND2_X1 U14550 ( .A1(n12786), .A2(n12785), .ZN(n12852) );
  NOR2_X1 U14551 ( .A1(n12852), .A2(n12910), .ZN(n12851) );
  AND2_X1 U14552 ( .A1(n12788), .A2(n12787), .ZN(n12793) );
  NAND2_X1 U14553 ( .A1(n12793), .A2(n12789), .ZN(n12790) );
  OAI21_X1 U14554 ( .B1(n12790), .B2(n12930), .A(n12805), .ZN(n12791) );
  NOR2_X1 U14555 ( .A1(n12792), .A2(n12791), .ZN(n12797) );
  INV_X1 U14556 ( .A(n12793), .ZN(n12794) );
  NAND3_X1 U14557 ( .A1(n12795), .A2(n9990), .A3(n12794), .ZN(n12796) );
  MUX2_X1 U14558 ( .A(n12797), .B(n12796), .S(n12910), .Z(n12803) );
  INV_X1 U14559 ( .A(n12800), .ZN(n12802) );
  NAND2_X1 U14560 ( .A1(n13483), .A2(n12798), .ZN(n12799) );
  AND2_X1 U14561 ( .A1(n12800), .A2(n12799), .ZN(n12801) );
  OAI22_X1 U14562 ( .A1(n12803), .A2(n12802), .B1(n12801), .B2(n12901), .ZN(
        n12804) );
  OAI211_X1 U14563 ( .C1(n12805), .C2(n12901), .A(n12804), .B(n7578), .ZN(
        n12808) );
  MUX2_X1 U14564 ( .A(n9647), .B(n12806), .S(n12910), .Z(n12807) );
  NAND3_X1 U14565 ( .A1(n12808), .A2(n12925), .A3(n12807), .ZN(n12813) );
  MUX2_X1 U14566 ( .A(n12810), .B(n12809), .S(n12901), .Z(n12811) );
  NAND3_X1 U14567 ( .A1(n12813), .A2(n12812), .A3(n12811), .ZN(n12818) );
  NAND2_X1 U14568 ( .A1(n13605), .A2(n12814), .ZN(n12815) );
  MUX2_X1 U14569 ( .A(n12816), .B(n12815), .S(n12910), .Z(n12817) );
  NAND3_X1 U14570 ( .A1(n12818), .A2(n12924), .A3(n12817), .ZN(n12822) );
  MUX2_X1 U14571 ( .A(n12820), .B(n12819), .S(n12901), .Z(n12821) );
  NAND3_X1 U14572 ( .A1(n12822), .A2(n12932), .A3(n12821), .ZN(n12827) );
  NAND2_X1 U14573 ( .A1(n13604), .A2(n12823), .ZN(n12824) );
  MUX2_X1 U14574 ( .A(n12825), .B(n12824), .S(n12910), .Z(n12826) );
  NAND3_X1 U14575 ( .A1(n12827), .A2(n7461), .A3(n12826), .ZN(n12831) );
  MUX2_X1 U14576 ( .A(n12829), .B(n7966), .S(n12910), .Z(n12830) );
  NAND2_X1 U14577 ( .A1(n12831), .A2(n12830), .ZN(n12838) );
  NAND2_X1 U14578 ( .A1(n12833), .A2(n12832), .ZN(n12835) );
  MUX2_X1 U14579 ( .A(n12835), .B(n12834), .S(n12910), .Z(n12836) );
  NAND2_X1 U14580 ( .A1(n12836), .A2(n12936), .ZN(n12837) );
  AOI21_X1 U14581 ( .B1(n12838), .B2(n12934), .A(n12837), .ZN(n12847) );
  NAND2_X1 U14582 ( .A1(n12844), .A2(n12839), .ZN(n12842) );
  NAND2_X1 U14583 ( .A1(n12843), .A2(n12840), .ZN(n12841) );
  MUX2_X1 U14584 ( .A(n12842), .B(n12841), .S(n12910), .Z(n12846) );
  MUX2_X1 U14585 ( .A(n12844), .B(n12843), .S(n12901), .Z(n12845) );
  OAI21_X1 U14586 ( .B1(n12847), .B2(n12846), .A(n12845), .ZN(n12850) );
  OR2_X1 U14587 ( .A1(n12848), .A2(n10012), .ZN(n12939) );
  INV_X1 U14588 ( .A(n12939), .ZN(n12849) );
  MUX2_X1 U14589 ( .A(n12851), .B(n12850), .S(n12849), .Z(n12854) );
  AND2_X1 U14590 ( .A1(n12852), .A2(n12910), .ZN(n12853) );
  OAI21_X1 U14591 ( .B1(n12854), .B2(n12853), .A(n13917), .ZN(n12858) );
  MUX2_X1 U14592 ( .A(n12856), .B(n12855), .S(n12910), .Z(n12857) );
  NAND3_X1 U14593 ( .A1(n12858), .A2(n13907), .A3(n12857), .ZN(n12859) );
  OAI21_X1 U14594 ( .B1(n12910), .B2(n12860), .A(n12859), .ZN(n12861) );
  NAND2_X1 U14595 ( .A1(n12861), .A2(n12942), .ZN(n12868) );
  INV_X1 U14596 ( .A(n12942), .ZN(n12863) );
  NOR2_X1 U14597 ( .A1(n12863), .A2(n12862), .ZN(n12866) );
  OAI211_X1 U14598 ( .C1(n7973), .C2(n12864), .A(n12874), .B(n12869), .ZN(
        n12865) );
  OAI21_X1 U14599 ( .B1(n12866), .B2(n12865), .A(n12910), .ZN(n12867) );
  NAND2_X1 U14600 ( .A1(n12868), .A2(n12867), .ZN(n12876) );
  NAND2_X1 U14601 ( .A1(n12876), .A2(n12871), .ZN(n12878) );
  INV_X1 U14602 ( .A(n12869), .ZN(n12873) );
  OAI211_X1 U14603 ( .C1(n12873), .C2(n12872), .A(n12871), .B(n12870), .ZN(
        n12875) );
  OAI21_X1 U14604 ( .B1(n12876), .B2(n12875), .A(n12874), .ZN(n12877) );
  MUX2_X1 U14605 ( .A(n12878), .B(n12877), .S(n12901), .Z(n12882) );
  MUX2_X1 U14606 ( .A(n12880), .B(n12879), .S(n12910), .Z(n12881) );
  OAI21_X1 U14607 ( .B1(n12882), .B2(n13852), .A(n12881), .ZN(n12883) );
  NAND2_X1 U14608 ( .A1(n12883), .A2(n7581), .ZN(n12888) );
  NOR2_X1 U14609 ( .A1(n14020), .A2(n13823), .ZN(n12885) );
  INV_X1 U14610 ( .A(n13401), .ZN(n12884) );
  MUX2_X1 U14611 ( .A(n12885), .B(n12884), .S(n12901), .Z(n12886) );
  INV_X1 U14612 ( .A(n12886), .ZN(n12887) );
  NAND3_X1 U14613 ( .A1(n12888), .A2(n13817), .A3(n12887), .ZN(n12892) );
  INV_X1 U14614 ( .A(n13808), .ZN(n12944) );
  NAND2_X1 U14615 ( .A1(n13833), .A2(n12901), .ZN(n12890) );
  NAND2_X1 U14616 ( .A1(n13806), .A2(n12910), .ZN(n12889) );
  MUX2_X1 U14617 ( .A(n12890), .B(n12889), .S(n14012), .Z(n12891) );
  NAND3_X1 U14618 ( .A1(n12892), .A2(n12944), .A3(n12891), .ZN(n12896) );
  NAND2_X1 U14619 ( .A1(n13811), .A2(n13824), .ZN(n12894) );
  MUX2_X1 U14620 ( .A(n12894), .B(n12893), .S(n12910), .Z(n12895) );
  NAND4_X1 U14621 ( .A1(n12897), .A2(n13791), .A3(n12896), .A4(n12895), .ZN(
        n12898) );
  INV_X1 U14622 ( .A(n12948), .ZN(n12903) );
  NAND3_X1 U14623 ( .A1(n13741), .A2(n13754), .A3(n12901), .ZN(n12902) );
  INV_X1 U14624 ( .A(n12904), .ZN(n12905) );
  OR2_X1 U14625 ( .A1(n12909), .A2(n12905), .ZN(n12912) );
  INV_X1 U14626 ( .A(n12906), .ZN(n12907) );
  AOI21_X1 U14627 ( .B1(n12909), .B2(n12908), .A(n12907), .ZN(n12911) );
  NAND2_X1 U14628 ( .A1(n13720), .A2(n12913), .ZN(n12949) );
  AND2_X1 U14629 ( .A1(n12915), .A2(n12914), .ZN(n12951) );
  INV_X1 U14630 ( .A(n12951), .ZN(n12916) );
  INV_X1 U14631 ( .A(n12955), .ZN(n12918) );
  INV_X1 U14632 ( .A(n12922), .ZN(n12923) );
  NAND4_X1 U14633 ( .A1(n7461), .A2(n12925), .A3(n12924), .A4(n12923), .ZN(
        n12929) );
  NAND3_X1 U14634 ( .A1(n12927), .A2(n7578), .A3(n12926), .ZN(n12928) );
  NOR2_X1 U14635 ( .A1(n12929), .A2(n12928), .ZN(n12935) );
  NOR2_X1 U14636 ( .A1(n12931), .A2(n12930), .ZN(n12933) );
  NAND4_X1 U14637 ( .A1(n12935), .A2(n12934), .A3(n12933), .A4(n12932), .ZN(
        n12938) );
  NAND2_X1 U14638 ( .A1(n13966), .A2(n12936), .ZN(n12937) );
  NOR4_X1 U14639 ( .A1(n12940), .A2(n12939), .A3(n12938), .A4(n12937), .ZN(
        n12941) );
  NAND4_X1 U14640 ( .A1(n13864), .A2(n13907), .A3(n12942), .A4(n12941), .ZN(
        n12943) );
  NOR3_X1 U14641 ( .A1(n13835), .A2(n13852), .A3(n12943), .ZN(n12945) );
  NAND4_X1 U14642 ( .A1(n13791), .A2(n12945), .A3(n12944), .A4(n13817), .ZN(
        n12946) );
  NOR4_X1 U14643 ( .A1(n12948), .A2(n13743), .A3(n12947), .A4(n12946), .ZN(
        n12950) );
  NAND4_X1 U14644 ( .A1(n12951), .A2(n12950), .A3(n12955), .A4(n12949), .ZN(
        n12952) );
  XNOR2_X1 U14645 ( .A(n12952), .B(n13694), .ZN(n12954) );
  NAND3_X1 U14646 ( .A1(n12961), .A2(n12960), .A3(n7429), .ZN(n12962) );
  OAI211_X1 U14647 ( .C1(n12963), .C2(n12965), .A(n12962), .B(P3_B_REG_SCAN_IN), .ZN(n12964) );
  INV_X1 U14648 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n12966) );
  NOR2_X1 U14649 ( .A1(n7428), .A2(n12966), .ZN(n12967) );
  INV_X1 U14650 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n12968) );
  NOR2_X1 U14651 ( .A1(n13284), .A2(n12968), .ZN(n12972) );
  INV_X1 U14652 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n15530) );
  NOR2_X1 U14653 ( .A1(n13256), .A2(n15530), .ZN(n12971) );
  INV_X1 U14654 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n12969) );
  NOR2_X1 U14655 ( .A1(n13279), .A2(n12969), .ZN(n12970) );
  OR3_X1 U14656 ( .A1(n12972), .A2(n12971), .A3(n12970), .ZN(n15531) );
  XNOR2_X1 U14657 ( .A(n15823), .B(n15531), .ZN(n13340) );
  OR2_X1 U14658 ( .A1(n13290), .A2(n15974), .ZN(n12974) );
  INV_X1 U14659 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n12978) );
  NAND2_X1 U14660 ( .A1(n13277), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n12977) );
  NAND2_X1 U14661 ( .A1(n13170), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n12976) );
  OAI211_X1 U14662 ( .C1(n13284), .C2(n12978), .A(n12977), .B(n12976), .ZN(
        n15586) );
  OAI21_X1 U14663 ( .B1(n15531), .B2(n12993), .A(n15586), .ZN(n12979) );
  INV_X1 U14664 ( .A(n12979), .ZN(n12989) );
  NAND2_X1 U14665 ( .A1(n12984), .A2(n13341), .ZN(n12981) );
  NAND2_X1 U14666 ( .A1(n12981), .A2(n12980), .ZN(n12982) );
  NAND2_X1 U14667 ( .A1(n12983), .A2(n12982), .ZN(n12988) );
  NAND2_X1 U14668 ( .A1(n12984), .A2(n15519), .ZN(n12985) );
  NAND2_X1 U14669 ( .A1(n12985), .A2(n16392), .ZN(n12986) );
  NAND2_X1 U14670 ( .A1(n15997), .A2(n12986), .ZN(n12987) );
  MUX2_X1 U14671 ( .A(n15526), .B(n12989), .S(n13105), .Z(n12990) );
  INV_X1 U14672 ( .A(n12990), .ZN(n13304) );
  OAI21_X1 U14673 ( .B1(n15531), .B2(n12999), .A(n15586), .ZN(n12991) );
  INV_X1 U14674 ( .A(n12991), .ZN(n12992) );
  MUX2_X1 U14675 ( .A(n12992), .B(n15526), .S(n13105), .Z(n13303) );
  NAND2_X1 U14676 ( .A1(n13304), .A2(n13303), .ZN(n13352) );
  INV_X1 U14677 ( .A(n13352), .ZN(n13000) );
  NAND2_X1 U14678 ( .A1(n12983), .A2(n12993), .ZN(n12994) );
  NAND2_X1 U14679 ( .A1(n12995), .A2(n12994), .ZN(n12997) );
  NAND2_X1 U14680 ( .A1(n12997), .A2(n12996), .ZN(n13360) );
  INV_X1 U14681 ( .A(n13360), .ZN(n13347) );
  NAND2_X1 U14682 ( .A1(n12999), .A2(n12998), .ZN(n13348) );
  INV_X1 U14683 ( .A(n13348), .ZN(n13358) );
  NAND2_X1 U14684 ( .A1(n15112), .A2(n13289), .ZN(n13002) );
  OR2_X1 U14685 ( .A1(n13290), .A2(n15977), .ZN(n13001) );
  NAND2_X1 U14686 ( .A1(n13170), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n13010) );
  INV_X1 U14687 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n13003) );
  OR2_X1 U14688 ( .A1(n13256), .A2(n13003), .ZN(n13009) );
  INV_X1 U14689 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n13121) );
  INV_X1 U14690 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13167) );
  INV_X1 U14691 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n15275) );
  NAND2_X1 U14692 ( .A1(n13209), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n13210) );
  NAND2_X1 U14693 ( .A1(n13245), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n13244) );
  NAND2_X1 U14694 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n13258), .ZN(n13257) );
  INV_X1 U14695 ( .A(n13257), .ZN(n13004) );
  NAND2_X1 U14696 ( .A1(n13004), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n13280) );
  INV_X1 U14697 ( .A(n13280), .ZN(n13005) );
  NAND2_X1 U14698 ( .A1(n13005), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n15588) );
  OR2_X1 U14699 ( .A1(n13282), .A2(n15588), .ZN(n13008) );
  INV_X1 U14700 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n13006) );
  OR2_X1 U14701 ( .A1(n13284), .A2(n13006), .ZN(n13007) );
  MUX2_X1 U14702 ( .A(n15830), .B(n15260), .S(n13105), .Z(n13297) );
  INV_X1 U14703 ( .A(n13297), .ZN(n13301) );
  NAND2_X1 U14704 ( .A1(n15118), .A2(n13289), .ZN(n13012) );
  OR2_X1 U14705 ( .A1(n7428), .A2(n15980), .ZN(n13011) );
  NAND2_X1 U14706 ( .A1(n13277), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n13020) );
  INV_X1 U14707 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n13013) );
  OR2_X1 U14708 ( .A1(n13279), .A2(n13013), .ZN(n13019) );
  INV_X1 U14709 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13014) );
  NAND2_X1 U14710 ( .A1(n13257), .A2(n13014), .ZN(n13015) );
  NAND2_X1 U14711 ( .A1(n13280), .A2(n13015), .ZN(n15618) );
  OR2_X1 U14712 ( .A1(n13282), .A2(n15618), .ZN(n13018) );
  INV_X1 U14713 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n13016) );
  OR2_X1 U14714 ( .A1(n13284), .A2(n13016), .ZN(n13017) );
  MUX2_X1 U14715 ( .A(n15840), .B(n15370), .S(n13105), .Z(n13275) );
  INV_X1 U14716 ( .A(n13275), .ZN(n13276) );
  NAND2_X1 U14717 ( .A1(n13021), .A2(n13345), .ZN(n13024) );
  NAND2_X1 U14718 ( .A1(n13022), .A2(n13105), .ZN(n13023) );
  NAND2_X1 U14719 ( .A1(n13024), .A2(n13023), .ZN(n13041) );
  OAI21_X1 U14720 ( .B1(n13310), .B2(n15384), .A(n13345), .ZN(n13037) );
  NAND2_X1 U14721 ( .A1(n8315), .A2(n13027), .ZN(n13032) );
  NAND2_X1 U14722 ( .A1(n15385), .A2(n13032), .ZN(n13029) );
  NAND2_X1 U14723 ( .A1(n13308), .A2(n13028), .ZN(n13031) );
  NAND3_X1 U14724 ( .A1(n13029), .A2(n7600), .A3(n13031), .ZN(n13030) );
  NAND2_X1 U14725 ( .A1(n13030), .A2(n7601), .ZN(n13035) );
  INV_X1 U14726 ( .A(n13031), .ZN(n13033) );
  OAI211_X1 U14727 ( .C1(n15385), .C2(n13033), .A(n13032), .B(n15384), .ZN(
        n13034) );
  NAND3_X1 U14728 ( .A1(n13035), .A2(n13105), .A3(n13034), .ZN(n13036) );
  OAI211_X1 U14729 ( .C1(n13038), .C2(n13037), .A(n13313), .B(n13036), .ZN(
        n13040) );
  NAND3_X1 U14730 ( .A1(n13041), .A2(n13040), .A3(n13039), .ZN(n13047) );
  NAND2_X1 U14731 ( .A1(n13042), .A2(n13105), .ZN(n13045) );
  NAND2_X1 U14732 ( .A1(n13043), .A2(n13345), .ZN(n13044) );
  AOI21_X1 U14733 ( .B1(n13045), .B2(n13044), .A(n13048), .ZN(n13046) );
  NAND3_X1 U14734 ( .A1(n13047), .A2(n13046), .A3(n13050), .ZN(n13052) );
  INV_X1 U14735 ( .A(n13048), .ZN(n13049) );
  MUX2_X1 U14736 ( .A(n13050), .B(n13049), .S(n13345), .Z(n13051) );
  NAND3_X1 U14737 ( .A1(n13052), .A2(n13051), .A3(n13311), .ZN(n13060) );
  OAI21_X1 U14738 ( .B1(n15380), .B2(n13345), .A(n13053), .ZN(n13057) );
  NAND2_X1 U14739 ( .A1(n15380), .A2(n13345), .ZN(n13055) );
  NAND2_X1 U14740 ( .A1(n13055), .A2(n13054), .ZN(n13056) );
  NAND2_X1 U14741 ( .A1(n13057), .A2(n13056), .ZN(n13058) );
  NAND3_X1 U14742 ( .A1(n13060), .A2(n13059), .A3(n13058), .ZN(n13064) );
  AND2_X1 U14743 ( .A1(n15379), .A2(n13105), .ZN(n13062) );
  OAI21_X1 U14744 ( .B1(n15379), .B2(n13105), .A(n16489), .ZN(n13061) );
  OAI21_X1 U14745 ( .B1(n13062), .B2(n16489), .A(n13061), .ZN(n13063) );
  NAND2_X1 U14746 ( .A1(n13064), .A2(n13063), .ZN(n13068) );
  MUX2_X1 U14747 ( .A(n15378), .B(n13065), .S(n13345), .Z(n13069) );
  NAND2_X1 U14748 ( .A1(n13068), .A2(n13069), .ZN(n13067) );
  MUX2_X1 U14749 ( .A(n15378), .B(n13065), .S(n13105), .Z(n13066) );
  NAND2_X1 U14750 ( .A1(n13067), .A2(n13066), .ZN(n13073) );
  INV_X1 U14751 ( .A(n13068), .ZN(n13071) );
  INV_X1 U14752 ( .A(n13069), .ZN(n13070) );
  NAND2_X1 U14753 ( .A1(n13071), .A2(n13070), .ZN(n13072) );
  NAND3_X1 U14754 ( .A1(n13073), .A2(n13072), .A3(n13320), .ZN(n13077) );
  AND2_X1 U14755 ( .A1(n15377), .A2(n13105), .ZN(n13075) );
  OAI21_X1 U14756 ( .B1(n15377), .B2(n13105), .A(n16526), .ZN(n13074) );
  OAI21_X1 U14757 ( .B1(n13075), .B2(n16526), .A(n13074), .ZN(n13076) );
  MUX2_X1 U14758 ( .A(n15376), .B(n13078), .S(n13345), .Z(n13080) );
  MUX2_X1 U14759 ( .A(n15376), .B(n13078), .S(n13105), .Z(n13079) );
  INV_X1 U14760 ( .A(n13080), .ZN(n13081) );
  MUX2_X1 U14761 ( .A(n15375), .B(n13082), .S(n13105), .Z(n13084) );
  MUX2_X1 U14762 ( .A(n15375), .B(n13082), .S(n13345), .Z(n13083) );
  INV_X1 U14763 ( .A(n13084), .ZN(n13085) );
  MUX2_X1 U14764 ( .A(n15374), .B(n13086), .S(n13345), .Z(n13088) );
  MUX2_X1 U14765 ( .A(n15374), .B(n13086), .S(n13105), .Z(n13087) );
  INV_X1 U14766 ( .A(n13088), .ZN(n13089) );
  MUX2_X1 U14767 ( .A(n15373), .B(n13090), .S(n13105), .Z(n13094) );
  NAND2_X1 U14768 ( .A1(n13093), .A2(n13094), .ZN(n13092) );
  MUX2_X1 U14769 ( .A(n15373), .B(n13090), .S(n13345), .Z(n13091) );
  NAND2_X1 U14770 ( .A1(n13092), .A2(n13091), .ZN(n13098) );
  INV_X1 U14771 ( .A(n13093), .ZN(n13096) );
  INV_X1 U14772 ( .A(n13094), .ZN(n13095) );
  NAND2_X1 U14773 ( .A1(n13096), .A2(n13095), .ZN(n13097) );
  MUX2_X1 U14774 ( .A(n15372), .B(n15940), .S(n13345), .Z(n13100) );
  MUX2_X1 U14775 ( .A(n15372), .B(n15940), .S(n13105), .Z(n13099) );
  INV_X1 U14776 ( .A(n13100), .ZN(n13101) );
  MUX2_X1 U14777 ( .A(n15371), .B(n13102), .S(n13105), .Z(n13104) );
  MUX2_X1 U14778 ( .A(n15371), .B(n13102), .S(n13345), .Z(n13103) );
  MUX2_X1 U14779 ( .A(n15540), .B(n15561), .S(n13345), .Z(n13107) );
  MUX2_X1 U14780 ( .A(n15540), .B(n15561), .S(n13105), .Z(n13106) );
  INV_X1 U14781 ( .A(n13107), .ZN(n13108) );
  NAND2_X1 U14782 ( .A1(n13109), .A2(n13289), .ZN(n13112) );
  AOI22_X1 U14783 ( .A1(n13155), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n13154), 
        .B2(n13110), .ZN(n13111) );
  MUX2_X1 U14784 ( .A(n15788), .B(n15919), .S(n13105), .Z(n13116) );
  NAND2_X1 U14785 ( .A1(n13115), .A2(n13116), .ZN(n13114) );
  MUX2_X1 U14786 ( .A(n15919), .B(n15788), .S(n13105), .Z(n13113) );
  NAND2_X1 U14787 ( .A1(n13114), .A2(n13113), .ZN(n13120) );
  INV_X1 U14788 ( .A(n13115), .ZN(n13118) );
  INV_X1 U14789 ( .A(n13116), .ZN(n13117) );
  NAND2_X1 U14790 ( .A1(n13118), .A2(n13117), .ZN(n13119) );
  AND2_X1 U14791 ( .A1(n13122), .A2(n13121), .ZN(n13123) );
  OR2_X1 U14792 ( .A1(n13123), .A2(n13138), .ZN(n15795) );
  AOI22_X1 U14793 ( .A1(n13170), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n13277), 
        .B2(P1_REG2_REG_17__SCAN_IN), .ZN(n13126) );
  OR2_X1 U14794 ( .A1(n13284), .A2(n13124), .ZN(n13125) );
  OAI211_X1 U14795 ( .C1(n15795), .C2(n13282), .A(n13126), .B(n13125), .ZN(
        n15768) );
  NAND2_X1 U14796 ( .A1(n13127), .A2(n13289), .ZN(n13131) );
  INV_X1 U14797 ( .A(n13128), .ZN(n13129) );
  AOI22_X1 U14798 ( .A1(n13155), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n13154), 
        .B2(n13129), .ZN(n13130) );
  MUX2_X1 U14799 ( .A(n15768), .B(n15909), .S(n13345), .Z(n13133) );
  MUX2_X1 U14800 ( .A(n15768), .B(n15909), .S(n13105), .Z(n13132) );
  INV_X1 U14801 ( .A(n13133), .ZN(n13134) );
  NAND2_X1 U14802 ( .A1(n13135), .A2(n13289), .ZN(n13137) );
  AOI22_X1 U14803 ( .A1(n13155), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n13154), 
        .B2(n15507), .ZN(n13136) );
  NOR2_X1 U14804 ( .A1(n13138), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13139) );
  OR2_X1 U14805 ( .A1(n13158), .A2(n13139), .ZN(n15775) );
  INV_X1 U14806 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n13142) );
  NAND2_X1 U14807 ( .A1(n13170), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n13141) );
  INV_X1 U14808 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15776) );
  OR2_X1 U14809 ( .A1(n13256), .A2(n15776), .ZN(n13140) );
  OAI211_X1 U14810 ( .C1(n13142), .C2(n13284), .A(n13141), .B(n13140), .ZN(
        n13143) );
  INV_X1 U14811 ( .A(n13143), .ZN(n13144) );
  OAI21_X1 U14812 ( .B1(n15775), .B2(n13282), .A(n13144), .ZN(n15790) );
  MUX2_X1 U14813 ( .A(n15778), .B(n15790), .S(n13345), .Z(n13148) );
  NAND2_X1 U14814 ( .A1(n13147), .A2(n13148), .ZN(n13146) );
  MUX2_X1 U14815 ( .A(n15778), .B(n15790), .S(n13105), .Z(n13145) );
  NAND2_X1 U14816 ( .A1(n13146), .A2(n13145), .ZN(n13152) );
  INV_X1 U14817 ( .A(n13147), .ZN(n13150) );
  INV_X1 U14818 ( .A(n13148), .ZN(n13149) );
  NAND2_X1 U14819 ( .A1(n13150), .A2(n13149), .ZN(n13151) );
  NAND2_X1 U14820 ( .A1(n13153), .A2(n13289), .ZN(n13157) );
  AOI22_X1 U14821 ( .A1(n13155), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n13341), 
        .B2(n13154), .ZN(n13156) );
  OR2_X1 U14822 ( .A1(n13158), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13159) );
  AND2_X1 U14823 ( .A1(n13168), .A2(n13159), .ZN(n15758) );
  INV_X1 U14824 ( .A(n13282), .ZN(n13212) );
  NAND2_X1 U14825 ( .A1(n15758), .A2(n13212), .ZN(n13164) );
  INV_X1 U14826 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n15505) );
  NAND2_X1 U14827 ( .A1(n13170), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n13161) );
  NAND2_X1 U14828 ( .A1(n13277), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n13160) );
  OAI211_X1 U14829 ( .C1(n15505), .C2(n13284), .A(n13161), .B(n13160), .ZN(
        n13162) );
  INV_X1 U14830 ( .A(n13162), .ZN(n13163) );
  NAND2_X1 U14831 ( .A1(n13164), .A2(n13163), .ZN(n15769) );
  MUX2_X1 U14832 ( .A(n15746), .B(n15769), .S(n13105), .Z(n13166) );
  MUX2_X1 U14833 ( .A(n15746), .B(n15769), .S(n13345), .Z(n13165) );
  NAND2_X1 U14834 ( .A1(n13168), .A2(n13167), .ZN(n13169) );
  AND2_X1 U14835 ( .A1(n13186), .A2(n13169), .ZN(n15740) );
  NAND2_X1 U14836 ( .A1(n15740), .A2(n13212), .ZN(n13175) );
  INV_X1 U14837 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n15895) );
  NAND2_X1 U14838 ( .A1(n13170), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n13172) );
  NAND2_X1 U14839 ( .A1(n13277), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n13171) );
  OAI211_X1 U14840 ( .C1(n15895), .C2(n13284), .A(n13172), .B(n13171), .ZN(
        n13173) );
  INV_X1 U14841 ( .A(n13173), .ZN(n13174) );
  NAND2_X1 U14842 ( .A1(n13175), .A2(n13174), .ZN(n15550) );
  NAND2_X1 U14843 ( .A1(n13176), .A2(n13289), .ZN(n13179) );
  OR2_X1 U14844 ( .A1(n13290), .A2(n13177), .ZN(n13178) );
  MUX2_X1 U14845 ( .A(n15550), .B(n15889), .S(n13105), .Z(n13181) );
  MUX2_X1 U14846 ( .A(n15550), .B(n15889), .S(n13345), .Z(n13180) );
  NAND2_X1 U14847 ( .A1(n13182), .A2(n13289), .ZN(n13185) );
  OR2_X1 U14848 ( .A1(n7428), .A2(n13183), .ZN(n13184) );
  AND2_X1 U14849 ( .A1(n13186), .A2(n15275), .ZN(n13187) );
  OR2_X1 U14850 ( .A1(n13187), .A2(n13196), .ZN(n15720) );
  INV_X1 U14851 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n13190) );
  NAND2_X1 U14852 ( .A1(n13170), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n13189) );
  NAND2_X1 U14853 ( .A1(n13277), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n13188) );
  OAI211_X1 U14854 ( .C1(n13190), .C2(n13284), .A(n13189), .B(n13188), .ZN(
        n13191) );
  INV_X1 U14855 ( .A(n13191), .ZN(n13192) );
  OAI21_X1 U14856 ( .B1(n15720), .B2(n13282), .A(n13192), .ZN(n15736) );
  MUX2_X1 U14857 ( .A(n15883), .B(n15736), .S(n13105), .Z(n13194) );
  MUX2_X1 U14858 ( .A(n15736), .B(n15883), .S(n13105), .Z(n13193) );
  INV_X1 U14859 ( .A(n13194), .ZN(n13195) );
  NOR2_X1 U14860 ( .A1(n13196), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n13197) );
  OR2_X1 U14861 ( .A1(n13209), .A2(n13197), .ZN(n15705) );
  INV_X1 U14862 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n13200) );
  NAND2_X1 U14863 ( .A1(n13170), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n13199) );
  NAND2_X1 U14864 ( .A1(n13277), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n13198) );
  OAI211_X1 U14865 ( .C1(n13200), .C2(n13284), .A(n13199), .B(n13198), .ZN(
        n13201) );
  INV_X1 U14866 ( .A(n13201), .ZN(n13202) );
  OAI21_X1 U14867 ( .B1(n15705), .B2(n13282), .A(n13202), .ZN(n15554) );
  MUX2_X1 U14868 ( .A(n15554), .B(n15698), .S(n13105), .Z(n13207) );
  MUX2_X1 U14869 ( .A(n15698), .B(n15554), .S(n13105), .Z(n13205) );
  INV_X1 U14870 ( .A(n13207), .ZN(n13208) );
  OR2_X1 U14871 ( .A1(n13209), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n13211) );
  AND2_X1 U14872 ( .A1(n13211), .A2(n13210), .ZN(n15684) );
  NAND2_X1 U14873 ( .A1(n15684), .A2(n13212), .ZN(n13217) );
  INV_X1 U14874 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n15873) );
  NAND2_X1 U14875 ( .A1(n13170), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n13214) );
  NAND2_X1 U14876 ( .A1(n13277), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n13213) );
  OAI211_X1 U14877 ( .C1(n15873), .C2(n13284), .A(n13214), .B(n13213), .ZN(
        n13215) );
  INV_X1 U14878 ( .A(n13215), .ZN(n13216) );
  NAND2_X1 U14879 ( .A1(n13217), .A2(n13216), .ZN(n15703) );
  NAND2_X1 U14880 ( .A1(n13218), .A2(n13289), .ZN(n13221) );
  OR2_X1 U14881 ( .A1(n7428), .A2(n13219), .ZN(n13220) );
  MUX2_X1 U14882 ( .A(n15703), .B(n15867), .S(n13345), .Z(n13225) );
  MUX2_X1 U14883 ( .A(n15703), .B(n15867), .S(n13105), .Z(n13222) );
  NAND2_X1 U14884 ( .A1(n13223), .A2(n13222), .ZN(n13229) );
  INV_X1 U14885 ( .A(n13224), .ZN(n13227) );
  INV_X1 U14886 ( .A(n13225), .ZN(n13226) );
  NAND2_X1 U14887 ( .A1(n13227), .A2(n13226), .ZN(n13228) );
  NAND2_X1 U14888 ( .A1(n13277), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n13237) );
  INV_X1 U14889 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n13230) );
  OR2_X1 U14890 ( .A1(n13279), .A2(n13230), .ZN(n13236) );
  OAI21_X1 U14891 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n13232), .A(n13231), 
        .ZN(n15670) );
  OR2_X1 U14892 ( .A1(n13282), .A2(n15670), .ZN(n13235) );
  INV_X1 U14893 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n13233) );
  OR2_X1 U14894 ( .A1(n13284), .A2(n13233), .ZN(n13234) );
  NAND4_X1 U14895 ( .A1(n13237), .A2(n13236), .A3(n13235), .A4(n13234), .ZN(
        n15577) );
  NAND2_X1 U14896 ( .A1(n15129), .A2(n13289), .ZN(n13239) );
  OR2_X1 U14897 ( .A1(n13290), .A2(n15993), .ZN(n13238) );
  MUX2_X1 U14898 ( .A(n15577), .B(n15859), .S(n13105), .Z(n13241) );
  MUX2_X1 U14899 ( .A(n15577), .B(n15859), .S(n13345), .Z(n13240) );
  INV_X1 U14900 ( .A(n13241), .ZN(n13242) );
  NAND2_X1 U14901 ( .A1(n13277), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n13250) );
  INV_X1 U14902 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n13243) );
  OR2_X1 U14903 ( .A1(n13284), .A2(n13243), .ZN(n13249) );
  OAI21_X1 U14904 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n13245), .A(n13244), 
        .ZN(n15656) );
  OR2_X1 U14905 ( .A1(n13282), .A2(n15656), .ZN(n13248) );
  INV_X1 U14906 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n13246) );
  OR2_X1 U14907 ( .A1(n13279), .A2(n13246), .ZN(n13247) );
  NAND4_X1 U14908 ( .A1(n13250), .A2(n13249), .A3(n13248), .A4(n13247), .ZN(
        n15667) );
  NAND2_X1 U14909 ( .A1(n15126), .A2(n13289), .ZN(n13252) );
  OR2_X1 U14910 ( .A1(n13290), .A2(n15988), .ZN(n13251) );
  MUX2_X1 U14911 ( .A(n15667), .B(n15853), .S(n13345), .Z(n13254) );
  MUX2_X1 U14912 ( .A(n15667), .B(n15853), .S(n13105), .Z(n13253) );
  INV_X1 U14913 ( .A(n13254), .ZN(n13255) );
  NAND2_X1 U14914 ( .A1(n13170), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n13263) );
  INV_X1 U14915 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n15643) );
  OR2_X1 U14916 ( .A1(n13256), .A2(n15643), .ZN(n13262) );
  OAI21_X1 U14917 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n13258), .A(n13257), 
        .ZN(n15639) );
  OR2_X1 U14918 ( .A1(n13282), .A2(n15639), .ZN(n13261) );
  INV_X1 U14919 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n13259) );
  OR2_X1 U14920 ( .A1(n13284), .A2(n13259), .ZN(n13260) );
  NAND4_X1 U14921 ( .A1(n13263), .A2(n13262), .A3(n13261), .A4(n13260), .ZN(
        n15614) );
  NAND2_X1 U14922 ( .A1(n15122), .A2(n13289), .ZN(n13265) );
  OR2_X1 U14923 ( .A1(n13290), .A2(n15983), .ZN(n13264) );
  MUX2_X1 U14924 ( .A(n15614), .B(n15847), .S(n13105), .Z(n13269) );
  NAND2_X1 U14925 ( .A1(n13268), .A2(n13269), .ZN(n13267) );
  MUX2_X1 U14926 ( .A(n15614), .B(n15847), .S(n13345), .Z(n13266) );
  NAND2_X1 U14927 ( .A1(n13267), .A2(n13266), .ZN(n13273) );
  INV_X1 U14928 ( .A(n13268), .ZN(n13271) );
  INV_X1 U14929 ( .A(n13269), .ZN(n13270) );
  NAND2_X1 U14930 ( .A1(n13271), .A2(n13270), .ZN(n13272) );
  MUX2_X1 U14931 ( .A(n15636), .B(n15621), .S(n13105), .Z(n13274) );
  NAND2_X1 U14932 ( .A1(n13277), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n13288) );
  INV_X1 U14933 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n13278) );
  OR2_X1 U14934 ( .A1(n13279), .A2(n13278), .ZN(n13287) );
  INV_X1 U14935 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n15263) );
  NAND2_X1 U14936 ( .A1(n13280), .A2(n15263), .ZN(n13281) );
  NAND2_X1 U14937 ( .A1(n15588), .A2(n13281), .ZN(n15603) );
  OR2_X1 U14938 ( .A1(n13282), .A2(n15603), .ZN(n13286) );
  INV_X1 U14939 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n13283) );
  OR2_X1 U14940 ( .A1(n13284), .A2(n13283), .ZN(n13285) );
  NAND4_X1 U14941 ( .A1(n13288), .A2(n13287), .A3(n13286), .A4(n13285), .ZN(
        n15613) );
  NAND2_X1 U14942 ( .A1(n13371), .A2(n13289), .ZN(n13292) );
  OR2_X1 U14943 ( .A1(n7428), .A2(n13372), .ZN(n13291) );
  MUX2_X1 U14944 ( .A(n15613), .B(n15837), .S(n13105), .Z(n13295) );
  INV_X1 U14945 ( .A(n13295), .ZN(n13294) );
  MUX2_X1 U14946 ( .A(n15837), .B(n15613), .S(n13105), .Z(n13293) );
  INV_X1 U14947 ( .A(n13298), .ZN(n13300) );
  INV_X1 U14948 ( .A(n15260), .ZN(n15369) );
  MUX2_X1 U14949 ( .A(n15369), .B(n13305), .S(n13105), .Z(n13296) );
  OAI21_X1 U14950 ( .B1(n13301), .B2(n13300), .A(n13299), .ZN(n13302) );
  INV_X1 U14951 ( .A(n13363), .ZN(n13365) );
  XNOR2_X1 U14952 ( .A(n13305), .B(n15260), .ZN(n15582) );
  XNOR2_X1 U14953 ( .A(n15526), .B(n15586), .ZN(n13338) );
  XNOR2_X1 U14954 ( .A(n15847), .B(n15653), .ZN(n15630) );
  XNOR2_X1 U14955 ( .A(n15853), .B(n15667), .ZN(n15650) );
  NAND2_X1 U14956 ( .A1(n15876), .A2(n15554), .ZN(n13306) );
  NAND2_X1 U14957 ( .A1(n15576), .A2(n13306), .ZN(n15575) );
  XNOR2_X1 U14958 ( .A(n15883), .B(n15736), .ZN(n15726) );
  NAND2_X1 U14959 ( .A1(n15905), .A2(n15790), .ZN(n15569) );
  INV_X1 U14960 ( .A(n15790), .ZN(n15753) );
  NAND2_X1 U14961 ( .A1(n15778), .A2(n15753), .ZN(n13307) );
  NAND2_X1 U14962 ( .A1(n15569), .A2(n13307), .ZN(n15764) );
  INV_X1 U14963 ( .A(n15768), .ZN(n15807) );
  XNOR2_X1 U14964 ( .A(n15909), .B(n15807), .ZN(n15785) );
  XNOR2_X1 U14965 ( .A(n15919), .B(n15788), .ZN(n15542) );
  NAND2_X1 U14966 ( .A1(n15385), .A2(n13308), .ZN(n13309) );
  NAND2_X1 U14967 ( .A1(n13310), .A2(n13309), .ZN(n16398) );
  NOR2_X1 U14968 ( .A1(n11122), .A2(n16398), .ZN(n13314) );
  NAND4_X1 U14969 ( .A1(n13314), .A2(n13313), .A3(n13312), .A4(n13311), .ZN(
        n13316) );
  NOR2_X1 U14970 ( .A1(n13316), .A2(n13315), .ZN(n13319) );
  NAND4_X1 U14971 ( .A1(n13320), .A2(n13319), .A3(n13318), .A4(n13317), .ZN(
        n13321) );
  NOR2_X1 U14972 ( .A1(n13322), .A2(n13321), .ZN(n13325) );
  NAND4_X1 U14973 ( .A1(n13326), .A2(n13325), .A3(n13324), .A4(n13323), .ZN(
        n13327) );
  NOR2_X1 U14974 ( .A1(n13328), .A2(n13327), .ZN(n13330) );
  NAND4_X1 U14975 ( .A1(n15542), .A2(n13330), .A3(n15559), .A4(n13329), .ZN(
        n13331) );
  NOR3_X1 U14976 ( .A1(n15764), .A2(n15785), .A3(n13331), .ZN(n13332) );
  XNOR2_X1 U14977 ( .A(n15889), .B(n15550), .ZN(n15741) );
  XNOR2_X1 U14978 ( .A(n15746), .B(n15769), .ZN(n15547) );
  NAND4_X1 U14979 ( .A1(n15726), .A2(n13332), .A3(n15741), .A4(n15547), .ZN(
        n13333) );
  NOR2_X1 U14980 ( .A1(n15575), .A2(n13333), .ZN(n13334) );
  XNOR2_X1 U14981 ( .A(n15859), .B(n15577), .ZN(n15664) );
  XNOR2_X1 U14982 ( .A(n15867), .B(n15703), .ZN(n15687) );
  NAND4_X1 U14983 ( .A1(n15650), .A2(n13334), .A3(n15664), .A4(n15687), .ZN(
        n13335) );
  NOR2_X1 U14984 ( .A1(n15630), .A2(n13335), .ZN(n13337) );
  NAND2_X1 U14985 ( .A1(n15837), .A2(n15613), .ZN(n15558) );
  OR2_X1 U14986 ( .A1(n15837), .A2(n15613), .ZN(n13336) );
  NAND2_X1 U14987 ( .A1(n15558), .A2(n13336), .ZN(n15598) );
  NAND4_X1 U14988 ( .A1(n13338), .A2(n13337), .A3(n15624), .A4(n15598), .ZN(
        n13339) );
  NOR3_X1 U14989 ( .A1(n13340), .A2(n15582), .A3(n13339), .ZN(n13342) );
  XNOR2_X1 U14990 ( .A(n13342), .B(n13341), .ZN(n13357) );
  INV_X1 U14991 ( .A(n15823), .ZN(n15533) );
  NOR2_X1 U14992 ( .A1(n13360), .A2(n15531), .ZN(n13344) );
  INV_X1 U14993 ( .A(n15531), .ZN(n13343) );
  NAND2_X1 U14994 ( .A1(n13343), .A2(n13105), .ZN(n13350) );
  MUX2_X1 U14995 ( .A(n13360), .B(n13344), .S(n13350), .Z(n13355) );
  NAND2_X1 U14996 ( .A1(n13347), .A2(n15531), .ZN(n13346) );
  NAND2_X1 U14997 ( .A1(n13345), .A2(n15531), .ZN(n13351) );
  MUX2_X1 U14998 ( .A(n13347), .B(n13346), .S(n13351), .Z(n13349) );
  OAI21_X1 U14999 ( .B1(n15533), .B2(n13349), .A(n13348), .ZN(n13354) );
  NOR2_X1 U15000 ( .A1(n15823), .A2(n13350), .ZN(n13361) );
  NOR2_X1 U15001 ( .A1(n15533), .A2(n13351), .ZN(n13362) );
  NOR4_X1 U15002 ( .A1(n13361), .A2(n13362), .A3(n13352), .A4(n13360), .ZN(
        n13353) );
  AOI211_X1 U15003 ( .C1(n15533), .C2(n13355), .A(n13354), .B(n13353), .ZN(
        n13356) );
  AOI21_X1 U15004 ( .B1(n13358), .B2(n13357), .A(n13356), .ZN(n13359) );
  INV_X1 U15005 ( .A(n13359), .ZN(n13364) );
  NOR3_X1 U15006 ( .A1(n13366), .A2(n15982), .A3(n15805), .ZN(n13368) );
  OAI21_X1 U15007 ( .B1(n13369), .B2(n15997), .A(P1_B_REG_SCAN_IN), .ZN(n13367) );
  OAI22_X1 U15008 ( .A1(n13370), .A2(n13369), .B1(n13368), .B2(n13367), .ZN(
        P1_U3242) );
  INV_X1 U15009 ( .A(n13371), .ZN(n15116) );
  OAI222_X1 U15010 ( .A1(n13373), .A2(P1_U3086), .B1(n15990), .B2(n15116), 
        .C1(n13372), .C2(n15987), .ZN(P1_U3327) );
  XNOR2_X1 U15011 ( .A(n13835), .B(n13428), .ZN(n13405) );
  INV_X1 U15012 ( .A(n13374), .ZN(n13375) );
  NAND2_X1 U15013 ( .A1(n13375), .A2(n8429), .ZN(n13544) );
  NAND2_X1 U15014 ( .A1(n13377), .A2(n13376), .ZN(n13543) );
  XOR2_X1 U15015 ( .A(n13428), .B(n13949), .Z(n13379) );
  INV_X1 U15016 ( .A(n13379), .ZN(n13546) );
  AND2_X1 U15017 ( .A1(n13543), .A2(n13546), .ZN(n13378) );
  NAND2_X1 U15018 ( .A1(n13544), .A2(n13378), .ZN(n13545) );
  NAND2_X1 U15019 ( .A1(n13379), .A2(n13968), .ZN(n13380) );
  NAND2_X1 U15020 ( .A1(n13545), .A2(n13380), .ZN(n13462) );
  XNOR2_X1 U15021 ( .A(n13469), .B(n13428), .ZN(n13381) );
  XNOR2_X1 U15022 ( .A(n13381), .B(n13550), .ZN(n13463) );
  OR2_X2 U15023 ( .A1(n13462), .A2(n13463), .ZN(n13460) );
  NAND2_X1 U15024 ( .A1(n13381), .A2(n13550), .ZN(n13382) );
  XNOR2_X1 U15025 ( .A(n13597), .B(n13428), .ZN(n13586) );
  XNOR2_X1 U15026 ( .A(n13912), .B(n13428), .ZN(n13508) );
  XNOR2_X1 U15027 ( .A(n13896), .B(n13428), .ZN(n13383) );
  XNOR2_X1 U15028 ( .A(n13383), .B(n13904), .ZN(n13519) );
  NAND2_X1 U15029 ( .A1(n13518), .A2(n13519), .ZN(n13386) );
  INV_X1 U15030 ( .A(n13383), .ZN(n13384) );
  NAND2_X1 U15031 ( .A1(n13384), .A2(n13904), .ZN(n13385) );
  NAND2_X1 U15032 ( .A1(n13386), .A2(n13385), .ZN(n13564) );
  XNOR2_X1 U15033 ( .A(n13884), .B(n13428), .ZN(n13387) );
  XNOR2_X1 U15034 ( .A(n13387), .B(n13868), .ZN(n13565) );
  NAND2_X1 U15035 ( .A1(n13564), .A2(n13565), .ZN(n13389) );
  NAND2_X1 U15036 ( .A1(n13387), .A2(n13892), .ZN(n13388) );
  XNOR2_X1 U15037 ( .A(n14027), .B(n13428), .ZN(n13390) );
  XNOR2_X1 U15038 ( .A(n13390), .B(n13856), .ZN(n13490) );
  XNOR2_X1 U15039 ( .A(n14023), .B(n13428), .ZN(n13391) );
  XNOR2_X1 U15040 ( .A(n13391), .B(n13867), .ZN(n13536) );
  INV_X1 U15041 ( .A(n13391), .ZN(n13392) );
  NAND2_X1 U15042 ( .A1(n13392), .A2(n13834), .ZN(n13393) );
  XOR2_X1 U15043 ( .A(n13405), .B(n13406), .Z(n13398) );
  AOI22_X1 U15044 ( .A1(n13834), .A2(n13589), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13395) );
  NAND2_X1 U15045 ( .A1(n13590), .A2(n13842), .ZN(n13394) );
  OAI211_X1 U15046 ( .C1(n13806), .C2(n13593), .A(n13395), .B(n13394), .ZN(
        n13396) );
  AOI21_X1 U15047 ( .B1(n14020), .B2(n13596), .A(n13396), .ZN(n13397) );
  OAI21_X1 U15048 ( .B1(n13398), .B2(n13599), .A(n13397), .ZN(P3_U3163) );
  INV_X1 U15049 ( .A(SI_27_), .ZN(n13399) );
  OAI222_X1 U15050 ( .A1(n14154), .A2(n13400), .B1(n14150), .B2(n13399), .C1(
        P3_U3151), .C2(n13671), .ZN(P3_U3268) );
  MUX2_X1 U15051 ( .A(n13402), .B(n13401), .S(n13428), .Z(n13407) );
  OR2_X1 U15052 ( .A1(n7465), .A2(n13407), .ZN(n13403) );
  AND2_X1 U15053 ( .A1(n7465), .A2(n13407), .ZN(n13408) );
  NAND3_X1 U15054 ( .A1(n13554), .A2(n13555), .A3(n13806), .ZN(n13556) );
  NAND2_X1 U15055 ( .A1(n13556), .A2(n13554), .ZN(n13412) );
  INV_X1 U15056 ( .A(n13412), .ZN(n13410) );
  XNOR2_X1 U15057 ( .A(n13811), .B(n13428), .ZN(n13411) );
  INV_X1 U15058 ( .A(n13411), .ZN(n13409) );
  NAND2_X1 U15059 ( .A1(n13410), .A2(n13409), .ZN(n13413) );
  NAND2_X1 U15060 ( .A1(n13412), .A2(n13411), .ZN(n13526) );
  XNOR2_X1 U15061 ( .A(n13801), .B(n13428), .ZN(n13414) );
  NAND2_X1 U15062 ( .A1(n13414), .A2(n13807), .ZN(n13497) );
  INV_X1 U15063 ( .A(n13414), .ZN(n13415) );
  NAND2_X1 U15064 ( .A1(n13415), .A2(n13602), .ZN(n13416) );
  XNOR2_X1 U15065 ( .A(n13507), .B(n13425), .ZN(n13417) );
  NAND2_X1 U15066 ( .A1(n13417), .A2(n13531), .ZN(n13420) );
  INV_X1 U15067 ( .A(n13417), .ZN(n13418) );
  NAND2_X1 U15068 ( .A1(n13418), .A2(n13795), .ZN(n13419) );
  NAND2_X1 U15069 ( .A1(n13500), .A2(n13420), .ZN(n13574) );
  XNOR2_X1 U15070 ( .A(n14081), .B(n13428), .ZN(n13422) );
  NOR2_X1 U15071 ( .A1(n13422), .A2(n13421), .ZN(n13423) );
  AOI21_X1 U15072 ( .B1(n13422), .B2(n13421), .A(n13423), .ZN(n13575) );
  INV_X1 U15073 ( .A(n13423), .ZN(n13424) );
  XNOR2_X1 U15074 ( .A(n13759), .B(n13425), .ZN(n13426) );
  NOR2_X1 U15075 ( .A1(n13426), .A2(n13768), .ZN(n13427) );
  AOI21_X1 U15076 ( .B1(n13426), .B2(n13768), .A(n13427), .ZN(n13453) );
  XNOR2_X1 U15077 ( .A(n13743), .B(n13428), .ZN(n13429) );
  OAI22_X1 U15078 ( .A1(n13733), .A2(n13568), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13430), .ZN(n13433) );
  INV_X1 U15079 ( .A(n13431), .ZN(n13739) );
  OAI22_X1 U15080 ( .A1(n13734), .A2(n13593), .B1(n13739), .B2(n13448), .ZN(
        n13432) );
  AOI211_X1 U15081 ( .C1(n13741), .C2(n13596), .A(n13433), .B(n13432), .ZN(
        n13434) );
  OAI21_X1 U15082 ( .B1(n13435), .B2(n13599), .A(n13434), .ZN(P3_U3160) );
  INV_X1 U15083 ( .A(SI_30_), .ZN(n13438) );
  INV_X1 U15084 ( .A(n13436), .ZN(n13437) );
  XOR2_X1 U15085 ( .A(n13442), .B(n13441), .Z(n13443) );
  NAND2_X1 U15086 ( .A1(n13443), .A2(n13576), .ZN(n13452) );
  AOI21_X1 U15087 ( .B1(n13605), .B2(n13589), .A(n13444), .ZN(n13451) );
  AOI22_X1 U15088 ( .A1(n13566), .A2(n13604), .B1(n13596), .B2(n13445), .ZN(
        n13450) );
  INV_X1 U15089 ( .A(n13446), .ZN(n13447) );
  OR2_X1 U15090 ( .A1(n13448), .A2(n13447), .ZN(n13449) );
  NAND4_X1 U15091 ( .A1(n13452), .A2(n13451), .A3(n13450), .A4(n13449), .ZN(
        P3_U3153) );
  NAND2_X1 U15092 ( .A1(n13454), .A2(n13576), .ZN(n13459) );
  INV_X1 U15093 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n13455) );
  OAI22_X1 U15094 ( .A1(n13779), .A2(n13568), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13455), .ZN(n13457) );
  NOR2_X1 U15095 ( .A1(n13754), .A2(n13593), .ZN(n13456) );
  AOI211_X1 U15096 ( .C1(n13758), .C2(n13590), .A(n13457), .B(n13456), .ZN(
        n13458) );
  OAI211_X1 U15097 ( .C1(n14076), .C2(n13582), .A(n13459), .B(n13458), .ZN(
        P3_U3154) );
  INV_X1 U15098 ( .A(n13460), .ZN(n13461) );
  AOI21_X1 U15099 ( .B1(n13463), .B2(n13462), .A(n13461), .ZN(n13471) );
  NAND2_X1 U15100 ( .A1(n13590), .A2(n13937), .ZN(n13466) );
  AOI21_X1 U15101 ( .B1(n13566), .B2(n13934), .A(n13464), .ZN(n13465) );
  OAI211_X1 U15102 ( .C1(n13467), .C2(n13568), .A(n13466), .B(n13465), .ZN(
        n13468) );
  AOI21_X1 U15103 ( .B1(n13469), .B2(n13596), .A(n13468), .ZN(n13470) );
  OAI21_X1 U15104 ( .B1(n13471), .B2(n13599), .A(n13470), .ZN(P3_U3155) );
  AOI21_X1 U15105 ( .B1(n13794), .B2(n13472), .A(n7441), .ZN(n13477) );
  AOI22_X1 U15106 ( .A1(n13833), .A2(n13589), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13474) );
  NAND2_X1 U15107 ( .A1(n13590), .A2(n13812), .ZN(n13473) );
  OAI211_X1 U15108 ( .C1(n13807), .C2(n13593), .A(n13474), .B(n13473), .ZN(
        n13475) );
  AOI21_X1 U15109 ( .B1(n13811), .B2(n13596), .A(n13475), .ZN(n13476) );
  OAI21_X1 U15110 ( .B1(n13477), .B2(n13599), .A(n13476), .ZN(P3_U3156) );
  OAI21_X1 U15111 ( .B1(n13480), .B2(n13479), .A(n13478), .ZN(n13481) );
  NAND3_X1 U15112 ( .A1(n7727), .A2(n13576), .A3(n13481), .ZN(n13489) );
  AOI21_X1 U15113 ( .B1(n13483), .B2(n13589), .A(n13482), .ZN(n13488) );
  AOI22_X1 U15114 ( .A1(n13485), .A2(n13566), .B1(n13596), .B2(n13484), .ZN(
        n13487) );
  NAND2_X1 U15115 ( .A1(n13590), .A2(n14472), .ZN(n13486) );
  NAND4_X1 U15116 ( .A1(n13489), .A2(n13488), .A3(n13487), .A4(n13486), .ZN(
        P3_U3158) );
  XNOR2_X1 U15117 ( .A(n13491), .B(n13490), .ZN(n13496) );
  INV_X1 U15118 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n14470) );
  NOR2_X1 U15119 ( .A1(n14470), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13705) );
  AOI21_X1 U15120 ( .B1(n13834), .B2(n13566), .A(n13705), .ZN(n13493) );
  NAND2_X1 U15121 ( .A1(n13590), .A2(n13869), .ZN(n13492) );
  OAI211_X1 U15122 ( .C1(n13868), .C2(n13568), .A(n13493), .B(n13492), .ZN(
        n13494) );
  AOI21_X1 U15123 ( .B1(n14027), .B2(n13596), .A(n13494), .ZN(n13495) );
  OAI21_X1 U15124 ( .B1(n13496), .B2(n13599), .A(n13495), .ZN(P3_U3159) );
  INV_X1 U15125 ( .A(n13497), .ZN(n13499) );
  NOR3_X1 U15126 ( .A1(n7710), .A2(n13499), .A3(n13498), .ZN(n13502) );
  INV_X1 U15127 ( .A(n13500), .ZN(n13501) );
  OAI21_X1 U15128 ( .B1(n13502), .B2(n13501), .A(n13576), .ZN(n13506) );
  AOI22_X1 U15129 ( .A1(n13602), .A2(n13589), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13503) );
  OAI21_X1 U15130 ( .B1(n13779), .B2(n13593), .A(n13503), .ZN(n13504) );
  AOI21_X1 U15131 ( .B1(n13784), .B2(n13590), .A(n13504), .ZN(n13505) );
  OAI211_X1 U15132 ( .C1(n13507), .C2(n13582), .A(n13506), .B(n13505), .ZN(
        P3_U3165) );
  XNOR2_X1 U15133 ( .A(n13508), .B(n13594), .ZN(n13509) );
  XNOR2_X1 U15134 ( .A(n13510), .B(n13509), .ZN(n13517) );
  NOR2_X1 U15135 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13511), .ZN(n13615) );
  AOI21_X1 U15136 ( .B1(n13904), .B2(n13566), .A(n13615), .ZN(n13513) );
  NAND2_X1 U15137 ( .A1(n13590), .A2(n13909), .ZN(n13512) );
  OAI211_X1 U15138 ( .C1(n13514), .C2(n13568), .A(n13513), .B(n13512), .ZN(
        n13515) );
  AOI21_X1 U15139 ( .B1(n14039), .B2(n13596), .A(n13515), .ZN(n13516) );
  OAI21_X1 U15140 ( .B1(n13517), .B2(n13599), .A(n13516), .ZN(P3_U3166) );
  XNOR2_X1 U15141 ( .A(n13518), .B(n13519), .ZN(n13525) );
  NAND2_X1 U15142 ( .A1(n13590), .A2(n13897), .ZN(n13522) );
  INV_X1 U15143 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n13520) );
  NOR2_X1 U15144 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13520), .ZN(n13652) );
  AOI21_X1 U15145 ( .B1(n13566), .B2(n13892), .A(n13652), .ZN(n13521) );
  OAI211_X1 U15146 ( .C1(n13594), .C2(n13568), .A(n13522), .B(n13521), .ZN(
        n13523) );
  AOI21_X1 U15147 ( .B1(n13896), .B2(n13596), .A(n13523), .ZN(n13524) );
  OAI21_X1 U15148 ( .B1(n13525), .B2(n13599), .A(n13524), .ZN(P3_U3168) );
  INV_X1 U15149 ( .A(n13801), .ZN(n14091) );
  INV_X1 U15150 ( .A(n13526), .ZN(n13528) );
  NOR3_X1 U15151 ( .A1(n7441), .A2(n13528), .A3(n13527), .ZN(n13529) );
  OAI21_X1 U15152 ( .B1(n13529), .B2(n7710), .A(n13576), .ZN(n13535) );
  INV_X1 U15153 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n13530) );
  OAI22_X1 U15154 ( .A1(n13824), .A2(n13568), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13530), .ZN(n13533) );
  NOR2_X1 U15155 ( .A1(n13531), .A2(n13593), .ZN(n13532) );
  AOI211_X1 U15156 ( .C1(n13800), .C2(n13590), .A(n13533), .B(n13532), .ZN(
        n13534) );
  OAI211_X1 U15157 ( .C1(n14091), .C2(n13582), .A(n13535), .B(n13534), .ZN(
        P3_U3169) );
  XNOR2_X1 U15158 ( .A(n13537), .B(n13536), .ZN(n13542) );
  NAND2_X1 U15159 ( .A1(n13590), .A2(n13860), .ZN(n13539) );
  AOI22_X1 U15160 ( .A1(n13566), .A2(n13855), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13538) );
  OAI211_X1 U15161 ( .C1(n13879), .C2(n13568), .A(n13539), .B(n13538), .ZN(
        n13540) );
  AOI21_X1 U15162 ( .B1(n14023), .B2(n13596), .A(n13540), .ZN(n13541) );
  OAI21_X1 U15163 ( .B1(n13542), .B2(n13599), .A(n13541), .ZN(P3_U3173) );
  AND2_X1 U15164 ( .A1(n13544), .A2(n13543), .ZN(n13547) );
  OAI211_X1 U15165 ( .C1(n13547), .C2(n13546), .A(n13576), .B(n13545), .ZN(
        n13553) );
  AOI21_X1 U15166 ( .B1(n13953), .B2(n13589), .A(n13548), .ZN(n13549) );
  OAI21_X1 U15167 ( .B1(n13550), .B2(n13593), .A(n13549), .ZN(n13551) );
  AOI21_X1 U15168 ( .B1(n13945), .B2(n13590), .A(n13551), .ZN(n13552) );
  OAI211_X1 U15169 ( .C1(n13582), .C2(n14055), .A(n13553), .B(n13552), .ZN(
        P3_U3174) );
  NAND2_X1 U15170 ( .A1(n13555), .A2(n13554), .ZN(n13558) );
  INV_X1 U15171 ( .A(n13556), .ZN(n13557) );
  AOI21_X1 U15172 ( .B1(n13833), .B2(n13558), .A(n13557), .ZN(n13563) );
  AOI22_X1 U15173 ( .A1(n13855), .A2(n13589), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13560) );
  NAND2_X1 U15174 ( .A1(n13590), .A2(n13819), .ZN(n13559) );
  OAI211_X1 U15175 ( .C1(n13824), .C2(n13593), .A(n13560), .B(n13559), .ZN(
        n13561) );
  AOI21_X1 U15176 ( .B1(n14012), .B2(n13596), .A(n13561), .ZN(n13562) );
  OAI21_X1 U15177 ( .B1(n13563), .B2(n13599), .A(n13562), .ZN(P3_U3175) );
  XNOR2_X1 U15178 ( .A(n13564), .B(n13565), .ZN(n13572) );
  NAND2_X1 U15179 ( .A1(n13566), .A2(n13856), .ZN(n13567) );
  NAND2_X1 U15180 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13666)
         );
  OAI211_X1 U15181 ( .C1(n13881), .C2(n13568), .A(n13567), .B(n13666), .ZN(
        n13570) );
  NOR2_X1 U15182 ( .A1(n13884), .A2(n13582), .ZN(n13569) );
  AOI211_X1 U15183 ( .C1(n13882), .C2(n13590), .A(n13570), .B(n13569), .ZN(
        n13571) );
  OAI21_X1 U15184 ( .B1(n13572), .B2(n13599), .A(n13571), .ZN(P3_U3178) );
  OAI21_X1 U15185 ( .B1(n13575), .B2(n13574), .A(n13573), .ZN(n13577) );
  NAND2_X1 U15186 ( .A1(n13577), .A2(n13576), .ZN(n13581) );
  AOI22_X1 U15187 ( .A1(n13795), .A2(n13589), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13578) );
  OAI21_X1 U15188 ( .B1(n13733), .B2(n13593), .A(n13578), .ZN(n13579) );
  AOI21_X1 U15189 ( .B1(n13773), .B2(n13590), .A(n13579), .ZN(n13580) );
  OAI211_X1 U15190 ( .C1(n14081), .C2(n13582), .A(n13581), .B(n13580), .ZN(
        P3_U3180) );
  INV_X1 U15191 ( .A(n13583), .ZN(n13585) );
  NAND2_X1 U15192 ( .A1(n13585), .A2(n13584), .ZN(n13587) );
  XNOR2_X1 U15193 ( .A(n13587), .B(n13586), .ZN(n13600) );
  INV_X1 U15194 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n13588) );
  NOR2_X1 U15195 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13588), .ZN(n16380) );
  AOI21_X1 U15196 ( .B1(n13955), .B2(n13589), .A(n16380), .ZN(n13592) );
  NAND2_X1 U15197 ( .A1(n13590), .A2(n13923), .ZN(n13591) );
  OAI211_X1 U15198 ( .C1(n13594), .C2(n13593), .A(n13592), .B(n13591), .ZN(
        n13595) );
  AOI21_X1 U15199 ( .B1(n13597), .B2(n13596), .A(n13595), .ZN(n13598) );
  OAI21_X1 U15200 ( .B1(n13600), .B2(n13599), .A(n13598), .ZN(P3_U3181) );
  MUX2_X1 U15201 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n13601), .S(n11644), .Z(
        P3_U3522) );
  MUX2_X1 U15202 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13768), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15203 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n13795), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15204 ( .A(n13602), .B(P3_DATAO_REG_24__SCAN_IN), .S(n13606), .Z(
        P3_U3515) );
  MUX2_X1 U15205 ( .A(n13833), .B(P3_DATAO_REG_22__SCAN_IN), .S(n13606), .Z(
        P3_U3513) );
  MUX2_X1 U15206 ( .A(n13855), .B(P3_DATAO_REG_21__SCAN_IN), .S(n13606), .Z(
        P3_U3512) );
  MUX2_X1 U15207 ( .A(n13856), .B(P3_DATAO_REG_19__SCAN_IN), .S(n13606), .Z(
        P3_U3510) );
  MUX2_X1 U15208 ( .A(n13892), .B(P3_DATAO_REG_18__SCAN_IN), .S(n13606), .Z(
        P3_U3509) );
  MUX2_X1 U15209 ( .A(n13904), .B(P3_DATAO_REG_17__SCAN_IN), .S(n13606), .Z(
        P3_U3508) );
  MUX2_X1 U15210 ( .A(n13920), .B(P3_DATAO_REG_16__SCAN_IN), .S(n13606), .Z(
        P3_U3507) );
  MUX2_X1 U15211 ( .A(n13934), .B(P3_DATAO_REG_15__SCAN_IN), .S(n13606), .Z(
        P3_U3506) );
  MUX2_X1 U15212 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n13955), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15213 ( .A(n13968), .B(P3_DATAO_REG_13__SCAN_IN), .S(n13606), .Z(
        P3_U3504) );
  MUX2_X1 U15214 ( .A(n13953), .B(P3_DATAO_REG_12__SCAN_IN), .S(n13606), .Z(
        P3_U3503) );
  MUX2_X1 U15215 ( .A(n13603), .B(P3_DATAO_REG_9__SCAN_IN), .S(n13606), .Z(
        P3_U3500) );
  MUX2_X1 U15216 ( .A(n13604), .B(P3_DATAO_REG_8__SCAN_IN), .S(n13606), .Z(
        P3_U3499) );
  MUX2_X1 U15217 ( .A(n13605), .B(P3_DATAO_REG_6__SCAN_IN), .S(n13606), .Z(
        P3_U3497) );
  MUX2_X1 U15218 ( .A(n13607), .B(P3_DATAO_REG_3__SCAN_IN), .S(n13606), .Z(
        P3_U3494) );
  MUX2_X1 U15219 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n10734), .S(P3_U3897), .Z(
        P3_U3492) );
  NOR2_X1 U15220 ( .A1(n13632), .A2(n13610), .ZN(n13611) );
  INV_X1 U15221 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n16373) );
  NOR2_X1 U15222 ( .A1(n16373), .A2(n16372), .ZN(n16371) );
  NOR2_X1 U15223 ( .A1(n13611), .A2(n16371), .ZN(n13614) );
  NAND2_X1 U15224 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n13649), .ZN(n13612) );
  OAI21_X1 U15225 ( .B1(P3_REG1_REG_16__SCAN_IN), .B2(n13649), .A(n13612), 
        .ZN(n13613) );
  AOI21_X1 U15226 ( .B1(n13614), .B2(n13613), .A(n13642), .ZN(n13641) );
  INV_X1 U15227 ( .A(n13649), .ZN(n13627) );
  INV_X1 U15228 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n16326) );
  INV_X1 U15229 ( .A(n13615), .ZN(n13616) );
  OAI21_X1 U15230 ( .B1(n16364), .B2(n16326), .A(n13616), .ZN(n13626) );
  NAND2_X1 U15231 ( .A1(n7489), .A2(n13632), .ZN(n13620) );
  OAI21_X1 U15232 ( .B1(n7489), .B2(n13632), .A(n13620), .ZN(n16369) );
  MUX2_X1 U15233 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n7429), .Z(n16370) );
  INV_X1 U15234 ( .A(n13620), .ZN(n13621) );
  NOR2_X1 U15235 ( .A1(n16368), .A2(n13621), .ZN(n13623) );
  MUX2_X1 U15236 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n7429), .Z(n13644) );
  XNOR2_X1 U15237 ( .A(n13644), .B(n13649), .ZN(n13622) );
  NOR2_X1 U15238 ( .A1(n13623), .A2(n13622), .ZN(n13647) );
  AOI21_X1 U15239 ( .B1(n13623), .B2(n13622), .A(n13647), .ZN(n13624) );
  NOR2_X1 U15240 ( .A1(n13624), .A2(n16376), .ZN(n13625) );
  AOI211_X1 U15241 ( .C1(n13707), .C2(n13627), .A(n13626), .B(n13625), .ZN(
        n13640) );
  OAI21_X1 U15242 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n13631), .A(n13630), 
        .ZN(n13633) );
  NOR2_X1 U15243 ( .A1(n13632), .A2(n13633), .ZN(n13634) );
  NOR2_X1 U15244 ( .A1(n16363), .A2(n16362), .ZN(n16361) );
  NOR2_X1 U15245 ( .A1(n13634), .A2(n16361), .ZN(n13637) );
  NAND2_X1 U15246 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n13649), .ZN(n13635) );
  OAI21_X1 U15247 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n13649), .A(n13635), 
        .ZN(n13636) );
  NOR2_X1 U15248 ( .A1(n13637), .A2(n13636), .ZN(n13648) );
  AOI21_X1 U15249 ( .B1(n13637), .B2(n13636), .A(n13648), .ZN(n13638) );
  OR2_X1 U15250 ( .A1(n13638), .A2(n16382), .ZN(n13639) );
  OAI211_X1 U15251 ( .C1(n13641), .C2(n16374), .A(n13640), .B(n13639), .ZN(
        P3_U3198) );
  INV_X1 U15252 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n14037) );
  AOI21_X1 U15253 ( .B1(n14037), .B2(n13643), .A(n13663), .ZN(n13659) );
  NOR2_X1 U15254 ( .A1(n13644), .A2(n13649), .ZN(n13646) );
  MUX2_X1 U15255 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n7429), .Z(n13669) );
  XNOR2_X1 U15256 ( .A(n13669), .B(n13668), .ZN(n13645) );
  NOR2_X1 U15257 ( .A1(n13667), .A2(n16376), .ZN(n13657) );
  OAI21_X1 U15258 ( .B1(n13647), .B2(n13646), .A(n13645), .ZN(n13656) );
  XOR2_X1 U15259 ( .A(n13678), .B(n13668), .Z(n13650) );
  AOI21_X1 U15260 ( .B1(n16036), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n13652), 
        .ZN(n13653) );
  OAI21_X1 U15261 ( .B1(n16367), .B2(n13668), .A(n13653), .ZN(n13654) );
  AOI211_X1 U15262 ( .C1(n13657), .C2(n13656), .A(n13655), .B(n13654), .ZN(
        n13658) );
  OAI21_X1 U15263 ( .B1(n13659), .B2(n16374), .A(n13658), .ZN(P3_U3199) );
  NAND2_X1 U15264 ( .A1(n13680), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n13689) );
  OR2_X1 U15265 ( .A1(n13680), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n13661) );
  AND2_X1 U15266 ( .A1(n13689), .A2(n13661), .ZN(n13662) );
  OAI21_X1 U15267 ( .B1(n13663), .B2(n7469), .A(n13662), .ZN(n13690) );
  INV_X1 U15268 ( .A(n13690), .ZN(n13665) );
  NOR3_X1 U15269 ( .A1(n13663), .A2(n7469), .A3(n13662), .ZN(n13664) );
  NOR2_X1 U15270 ( .A1(n13665), .A2(n13664), .ZN(n13688) );
  INV_X1 U15271 ( .A(n13680), .ZN(n13677) );
  INV_X1 U15272 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n16345) );
  OAI21_X1 U15273 ( .B1(n16364), .B2(n16345), .A(n13666), .ZN(n13676) );
  NAND2_X1 U15274 ( .A1(n13670), .A2(n13677), .ZN(n13700) );
  OAI21_X1 U15275 ( .B1(n13670), .B2(n13677), .A(n13700), .ZN(n13673) );
  MUX2_X1 U15276 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n7429), .Z(n13672) );
  NOR2_X1 U15277 ( .A1(n13673), .A2(n13672), .ZN(n13702) );
  AOI21_X1 U15278 ( .B1(n13673), .B2(n13672), .A(n13702), .ZN(n13674) );
  NOR2_X1 U15279 ( .A1(n13674), .A2(n16376), .ZN(n13675) );
  AOI211_X1 U15280 ( .C1(n13707), .C2(n13677), .A(n13676), .B(n13675), .ZN(
        n13687) );
  NAND2_X1 U15281 ( .A1(n13680), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n13692) );
  OR2_X1 U15282 ( .A1(n13680), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n13681) );
  AND2_X1 U15283 ( .A1(n13692), .A2(n13681), .ZN(n13682) );
  OAI21_X1 U15284 ( .B1(n13683), .B2(n13679), .A(n13682), .ZN(n13693) );
  INV_X1 U15285 ( .A(n13693), .ZN(n13685) );
  NOR3_X1 U15286 ( .A1(n13683), .A2(n13679), .A3(n13682), .ZN(n13684) );
  OAI21_X1 U15287 ( .B1(n13685), .B2(n13684), .A(n13712), .ZN(n13686) );
  OAI211_X1 U15288 ( .C1(n13688), .C2(n16374), .A(n13687), .B(n13686), .ZN(
        P3_U3200) );
  NAND2_X1 U15289 ( .A1(n13690), .A2(n13689), .ZN(n13691) );
  XNOR2_X1 U15290 ( .A(n13694), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13699) );
  XNOR2_X1 U15291 ( .A(n13691), .B(n13699), .ZN(n13714) );
  NAND2_X1 U15292 ( .A1(n13693), .A2(n13692), .ZN(n13696) );
  XNOR2_X1 U15293 ( .A(n13694), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13698) );
  INV_X1 U15294 ( .A(n13698), .ZN(n13695) );
  MUX2_X1 U15295 ( .A(n13699), .B(n13698), .S(n13697), .Z(n13704) );
  INV_X1 U15296 ( .A(n13700), .ZN(n13701) );
  NOR2_X1 U15297 ( .A1(n13702), .A2(n13701), .ZN(n13703) );
  XOR2_X1 U15298 ( .A(n13704), .B(n13703), .Z(n13710) );
  AOI21_X1 U15299 ( .B1(n16036), .B2(P3_ADDR_REG_19__SCAN_IN), .A(n13705), 
        .ZN(n13709) );
  NAND2_X1 U15300 ( .A1(n13707), .A2(n13706), .ZN(n13708) );
  OAI211_X1 U15301 ( .C1(n13710), .C2(n16376), .A(n13709), .B(n13708), .ZN(
        n13711) );
  OAI21_X1 U15302 ( .B1(n13714), .B2(n16374), .A(n13713), .ZN(P3_U3201) );
  NOR2_X1 U15303 ( .A1(n13717), .A2(n13716), .ZN(n14065) );
  NOR2_X1 U15304 ( .A1(n13718), .A2(n13946), .ZN(n13725) );
  NOR3_X1 U15305 ( .A1(n14065), .A2(n13958), .A3(n13725), .ZN(n13722) );
  NOR2_X1 U15306 ( .A1(n13977), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13719) );
  OAI22_X1 U15307 ( .A1(n14067), .A2(n13940), .B1(n13722), .B2(n13719), .ZN(
        P3_U3202) );
  NOR2_X1 U15308 ( .A1(n13977), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13721) );
  OAI22_X1 U15309 ( .A1(n14070), .A2(n13940), .B1(n13722), .B2(n13721), .ZN(
        P3_U3203) );
  INV_X1 U15310 ( .A(n13723), .ZN(n13730) );
  AOI21_X1 U15311 ( .B1(n13910), .B2(P3_REG2_REG_29__SCAN_IN), .A(n13725), 
        .ZN(n13726) );
  OAI21_X1 U15312 ( .B1(n13727), .B2(n13940), .A(n13726), .ZN(n13728) );
  AOI21_X1 U15313 ( .B1(n13724), .B2(n13977), .A(n13728), .ZN(n13729) );
  OAI21_X1 U15314 ( .B1(n13730), .B2(n13963), .A(n13729), .ZN(P3_U3204) );
  OAI211_X1 U15315 ( .C1(n13732), .C2(n13743), .A(n13731), .B(n13973), .ZN(
        n13737) );
  OAI22_X1 U15316 ( .A1(n13734), .A2(n13880), .B1(n13733), .B2(n13970), .ZN(
        n13735) );
  INV_X1 U15317 ( .A(n13735), .ZN(n13736) );
  OAI22_X1 U15318 ( .A1(n13739), .A2(n13946), .B1(n13977), .B2(n13738), .ZN(
        n13740) );
  AOI21_X1 U15319 ( .B1(n13741), .B2(n13981), .A(n13740), .ZN(n13745) );
  XNOR2_X1 U15320 ( .A(n13742), .B(n13743), .ZN(n13988) );
  NAND2_X1 U15321 ( .A1(n13988), .A2(n13942), .ZN(n13744) );
  OAI211_X1 U15322 ( .C1(n13990), .C2(n13958), .A(n13745), .B(n13744), .ZN(
        P3_U3205) );
  XNOR2_X1 U15323 ( .A(n13746), .B(n13750), .ZN(n13747) );
  NAND2_X1 U15324 ( .A1(n13751), .A2(n13750), .ZN(n13752) );
  NAND2_X1 U15325 ( .A1(n13749), .A2(n13752), .ZN(n13753) );
  NAND2_X1 U15326 ( .A1(n13753), .A2(n13973), .ZN(n13757) );
  OAI22_X1 U15327 ( .A1(n13754), .A2(n13880), .B1(n13779), .B2(n13970), .ZN(
        n13755) );
  INV_X1 U15328 ( .A(n13755), .ZN(n13756) );
  OAI211_X1 U15329 ( .C1(n14015), .C2(n13747), .A(n13757), .B(n13756), .ZN(
        n14075) );
  MUX2_X1 U15330 ( .A(n14075), .B(P3_REG2_REG_27__SCAN_IN), .S(n13910), .Z(
        n13762) );
  AOI22_X1 U15331 ( .A1(n13759), .A2(n13981), .B1(n13980), .B2(n13758), .ZN(
        n13760) );
  OAI21_X1 U15332 ( .B1(n13747), .B2(n13984), .A(n13760), .ZN(n13761) );
  INV_X1 U15333 ( .A(n14083), .ZN(n13999) );
  INV_X1 U15334 ( .A(n13764), .ZN(n13765) );
  XNOR2_X1 U15335 ( .A(n13766), .B(n13765), .ZN(n13767) );
  NAND2_X1 U15336 ( .A1(n13767), .A2(n13973), .ZN(n13771) );
  AOI22_X1 U15337 ( .A1(n13768), .A2(n13967), .B1(n13954), .B2(n13795), .ZN(
        n13770) );
  NAND2_X1 U15338 ( .A1(n14083), .A2(n14052), .ZN(n13769) );
  MUX2_X1 U15339 ( .A(n14079), .B(n13772), .S(n13910), .Z(n13775) );
  AOI22_X1 U15340 ( .A1(n13996), .A2(n13981), .B1(n13980), .B2(n13773), .ZN(
        n13774) );
  OAI211_X1 U15341 ( .C1(n13999), .C2(n13984), .A(n13775), .B(n13774), .ZN(
        P3_U3207) );
  AOI21_X1 U15342 ( .B1(n13778), .B2(n13777), .A(n13878), .ZN(n13782) );
  OAI22_X1 U15343 ( .A1(n13779), .A2(n13880), .B1(n13807), .B2(n13970), .ZN(
        n13780) );
  AOI21_X1 U15344 ( .B1(n13782), .B2(n13781), .A(n13780), .ZN(n13783) );
  OAI21_X1 U15345 ( .B1(n14015), .B2(n14089), .A(n13783), .ZN(n14000) );
  NAND2_X1 U15346 ( .A1(n14000), .A2(n13977), .ZN(n13789) );
  INV_X1 U15347 ( .A(n13784), .ZN(n13786) );
  OAI22_X1 U15348 ( .A1(n13786), .A2(n13946), .B1(n13977), .B2(n13785), .ZN(
        n13787) );
  AOI21_X1 U15349 ( .B1(n14001), .B2(n13981), .A(n13787), .ZN(n13788) );
  OAI211_X1 U15350 ( .C1(n14089), .C2(n13984), .A(n13789), .B(n13788), .ZN(
        P3_U3208) );
  XNOR2_X1 U15351 ( .A(n13792), .B(n13791), .ZN(n13793) );
  NAND2_X1 U15352 ( .A1(n13793), .A2(n13973), .ZN(n13797) );
  AOI22_X1 U15353 ( .A1(n13795), .A2(n13967), .B1(n13954), .B2(n13794), .ZN(
        n13796) );
  OAI211_X1 U15354 ( .C1(n14015), .C2(n14092), .A(n13797), .B(n13796), .ZN(
        n14090) );
  INV_X1 U15355 ( .A(n14090), .ZN(n13799) );
  MUX2_X1 U15356 ( .A(n13799), .B(n13798), .S(n13910), .Z(n13803) );
  AOI22_X1 U15357 ( .A1(n13801), .A2(n13981), .B1(n13980), .B2(n13800), .ZN(
        n13802) );
  OAI211_X1 U15358 ( .C1(n14092), .C2(n13984), .A(n13803), .B(n13802), .ZN(
        P3_U3209) );
  XNOR2_X1 U15359 ( .A(n13804), .B(n13808), .ZN(n13805) );
  OAI222_X1 U15360 ( .A1(n13880), .A2(n13807), .B1(n13970), .B2(n13806), .C1(
        n13878), .C2(n13805), .ZN(n14007) );
  INV_X1 U15361 ( .A(n14008), .ZN(n13810) );
  AND2_X1 U15362 ( .A1(n13809), .A2(n13808), .ZN(n14006) );
  NOR3_X1 U15363 ( .A1(n13810), .A2(n14006), .A3(n13963), .ZN(n13815) );
  INV_X1 U15364 ( .A(n13811), .ZN(n14098) );
  AOI22_X1 U15365 ( .A1(n13958), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n13980), 
        .B2(n13812), .ZN(n13813) );
  OAI21_X1 U15366 ( .B1(n14098), .B2(n13940), .A(n13813), .ZN(n13814) );
  AOI211_X1 U15367 ( .C1(n14007), .C2(n13977), .A(n13815), .B(n13814), .ZN(
        n13816) );
  INV_X1 U15368 ( .A(n13816), .ZN(P3_U3210) );
  XNOR2_X1 U15369 ( .A(n13818), .B(n7982), .ZN(n14102) );
  INV_X1 U15370 ( .A(n13819), .ZN(n13820) );
  OAI22_X1 U15371 ( .A1(n13977), .A2(n13821), .B1(n13820), .B2(n13946), .ZN(
        n13828) );
  XNOR2_X1 U15372 ( .A(n13822), .B(n7982), .ZN(n13826) );
  OAI22_X1 U15373 ( .A1(n13824), .A2(n13880), .B1(n13823), .B2(n13970), .ZN(
        n13825) );
  AOI21_X1 U15374 ( .B1(n13826), .B2(n13973), .A(n13825), .ZN(n14014) );
  NOR2_X1 U15375 ( .A1(n14014), .A2(n13958), .ZN(n13827) );
  AOI211_X1 U15376 ( .C1(n13981), .C2(n14012), .A(n13828), .B(n13827), .ZN(
        n13829) );
  OAI21_X1 U15377 ( .B1(n14102), .B2(n13963), .A(n13829), .ZN(P3_U3211) );
  NAND2_X1 U15378 ( .A1(n13853), .A2(n13852), .ZN(n13831) );
  NAND2_X1 U15379 ( .A1(n13831), .A2(n13830), .ZN(n13832) );
  XNOR2_X1 U15380 ( .A(n13832), .B(n13835), .ZN(n13841) );
  AOI22_X1 U15381 ( .A1(n13834), .A2(n13954), .B1(n13967), .B2(n13833), .ZN(
        n13840) );
  NAND2_X1 U15382 ( .A1(n13836), .A2(n13835), .ZN(n13837) );
  NAND2_X1 U15383 ( .A1(n13838), .A2(n13837), .ZN(n14018) );
  NAND2_X1 U15384 ( .A1(n14018), .A2(n14052), .ZN(n13839) );
  OAI211_X1 U15385 ( .C1(n13841), .C2(n13878), .A(n13840), .B(n13839), .ZN(
        n14019) );
  INV_X1 U15386 ( .A(n14019), .ZN(n13848) );
  INV_X1 U15387 ( .A(n14020), .ZN(n13844) );
  AOI22_X1 U15388 ( .A1(n13958), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n13980), 
        .B2(n13842), .ZN(n13843) );
  OAI21_X1 U15389 ( .B1(n13844), .B2(n13940), .A(n13843), .ZN(n13845) );
  AOI21_X1 U15390 ( .B1(n14018), .B2(n13846), .A(n13845), .ZN(n13847) );
  OAI21_X1 U15391 ( .B1(n13848), .B2(n13958), .A(n13847), .ZN(P3_U3212) );
  NAND2_X1 U15392 ( .A1(n13849), .A2(n13852), .ZN(n13850) );
  NAND2_X1 U15393 ( .A1(n13851), .A2(n13850), .ZN(n14110) );
  XNOR2_X1 U15394 ( .A(n13853), .B(n7579), .ZN(n13854) );
  NAND2_X1 U15395 ( .A1(n13854), .A2(n13973), .ZN(n13858) );
  AOI22_X1 U15396 ( .A1(n13954), .A2(n13856), .B1(n13855), .B2(n13967), .ZN(
        n13857) );
  OAI211_X1 U15397 ( .C1(n14015), .C2(n14110), .A(n13858), .B(n13857), .ZN(
        n14107) );
  MUX2_X1 U15398 ( .A(P3_REG2_REG_20__SCAN_IN), .B(n14107), .S(n13977), .Z(
        n13859) );
  INV_X1 U15399 ( .A(n13859), .ZN(n13862) );
  AOI22_X1 U15400 ( .A1(n14023), .A2(n13981), .B1(n13980), .B2(n13860), .ZN(
        n13861) );
  OAI211_X1 U15401 ( .C1(n14110), .C2(n13984), .A(n13862), .B(n13861), .ZN(
        P3_U3213) );
  XOR2_X1 U15402 ( .A(n13863), .B(n13864), .Z(n14029) );
  XNOR2_X1 U15403 ( .A(n13865), .B(n13864), .ZN(n13866) );
  OAI222_X1 U15404 ( .A1(n13970), .A2(n13868), .B1(n13880), .B2(n13867), .C1(
        n13878), .C2(n13866), .ZN(n14026) );
  AOI22_X1 U15405 ( .A1(n13958), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n13980), 
        .B2(n13869), .ZN(n13870) );
  OAI21_X1 U15406 ( .B1(n13871), .B2(n13940), .A(n13870), .ZN(n13872) );
  AOI21_X1 U15407 ( .B1(n14026), .B2(n13977), .A(n13872), .ZN(n13873) );
  OAI21_X1 U15408 ( .B1(n13963), .B2(n14029), .A(n13873), .ZN(P3_U3214) );
  XOR2_X1 U15409 ( .A(n13874), .B(n13876), .Z(n14033) );
  AOI21_X1 U15410 ( .B1(n13876), .B2(n13875), .A(n10019), .ZN(n13877) );
  OAI222_X1 U15411 ( .A1(n13970), .A2(n13881), .B1(n13880), .B2(n13879), .C1(
        n13878), .C2(n13877), .ZN(n14030) );
  AOI22_X1 U15412 ( .A1(n13958), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n13980), 
        .B2(n13882), .ZN(n13883) );
  OAI21_X1 U15413 ( .B1(n13884), .B2(n13940), .A(n13883), .ZN(n13885) );
  AOI21_X1 U15414 ( .B1(n14030), .B2(n13977), .A(n13885), .ZN(n13886) );
  OAI21_X1 U15415 ( .B1(n13963), .B2(n14033), .A(n13886), .ZN(P3_U3215) );
  XNOR2_X1 U15416 ( .A(n13888), .B(n13887), .ZN(n14036) );
  INV_X1 U15417 ( .A(n14036), .ZN(n13901) );
  NAND2_X1 U15418 ( .A1(n13889), .A2(n13973), .ZN(n13895) );
  AOI21_X1 U15419 ( .B1(n13902), .B2(n13891), .A(n13890), .ZN(n13894) );
  AOI22_X1 U15420 ( .A1(n13967), .A2(n13892), .B1(n13920), .B2(n13954), .ZN(
        n13893) );
  OAI21_X1 U15421 ( .B1(n13895), .B2(n13894), .A(n13893), .ZN(n14035) );
  INV_X1 U15422 ( .A(n13896), .ZN(n14118) );
  AOI22_X1 U15423 ( .A1(n13958), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n13980), 
        .B2(n13897), .ZN(n13898) );
  OAI21_X1 U15424 ( .B1(n14118), .B2(n13940), .A(n13898), .ZN(n13899) );
  AOI21_X1 U15425 ( .B1(n14035), .B2(n13977), .A(n13899), .ZN(n13900) );
  OAI21_X1 U15426 ( .B1(n13963), .B2(n13901), .A(n13900), .ZN(P3_U3216) );
  OAI21_X1 U15427 ( .B1(n13903), .B2(n10016), .A(n13902), .ZN(n13905) );
  AOI222_X1 U15428 ( .A1(n13973), .A2(n13905), .B1(n13934), .B2(n13954), .C1(
        n13904), .C2(n13967), .ZN(n14043) );
  OAI21_X1 U15429 ( .B1(n13908), .B2(n13907), .A(n13906), .ZN(n14041) );
  AOI22_X1 U15430 ( .A1(n13910), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n13980), 
        .B2(n13909), .ZN(n13911) );
  OAI21_X1 U15431 ( .B1(n13912), .B2(n13940), .A(n13911), .ZN(n13913) );
  AOI21_X1 U15432 ( .B1(n14041), .B2(n13942), .A(n13913), .ZN(n13914) );
  OAI21_X1 U15433 ( .B1(n14043), .B2(n13958), .A(n13914), .ZN(P3_U3217) );
  XNOR2_X1 U15434 ( .A(n13915), .B(n13917), .ZN(n14045) );
  INV_X1 U15435 ( .A(n14045), .ZN(n13927) );
  NAND3_X1 U15436 ( .A1(n13933), .A2(n13917), .A3(n13916), .ZN(n13918) );
  NAND3_X1 U15437 ( .A1(n13919), .A2(n13973), .A3(n13918), .ZN(n13922) );
  AOI22_X1 U15438 ( .A1(n13955), .A2(n13954), .B1(n13967), .B2(n13920), .ZN(
        n13921) );
  NAND2_X1 U15439 ( .A1(n13922), .A2(n13921), .ZN(n14044) );
  AOI22_X1 U15440 ( .A1(n13958), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n13980), 
        .B2(n13923), .ZN(n13924) );
  OAI21_X1 U15441 ( .B1(n14123), .B2(n13940), .A(n13924), .ZN(n13925) );
  AOI21_X1 U15442 ( .B1(n14044), .B2(n13977), .A(n13925), .ZN(n13926) );
  OAI21_X1 U15443 ( .B1(n13963), .B2(n13927), .A(n13926), .ZN(P3_U3218) );
  XNOR2_X1 U15444 ( .A(n13928), .B(n13931), .ZN(n14048) );
  NAND3_X1 U15445 ( .A1(n13952), .A2(n13931), .A3(n13930), .ZN(n13932) );
  NAND3_X1 U15446 ( .A1(n13933), .A2(n13973), .A3(n13932), .ZN(n13936) );
  AOI22_X1 U15447 ( .A1(n13967), .A2(n13934), .B1(n13968), .B2(n13954), .ZN(
        n13935) );
  NAND2_X1 U15448 ( .A1(n13936), .A2(n13935), .ZN(n14047) );
  NAND2_X1 U15449 ( .A1(n14047), .A2(n13977), .ZN(n13939) );
  AOI22_X1 U15450 ( .A1(n13958), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n13980), 
        .B2(n13937), .ZN(n13938) );
  OAI211_X1 U15451 ( .C1(n13940), .C2(n14127), .A(n13939), .B(n13938), .ZN(
        n13941) );
  AOI21_X1 U15452 ( .B1(n13942), .B2(n14048), .A(n13941), .ZN(n13943) );
  INV_X1 U15453 ( .A(n13943), .ZN(P3_U3219) );
  XNOR2_X1 U15454 ( .A(n13944), .B(n13949), .ZN(n14130) );
  INV_X1 U15455 ( .A(n14130), .ZN(n14058) );
  INV_X1 U15456 ( .A(n13945), .ZN(n13947) );
  OAI22_X1 U15457 ( .A1(n13977), .A2(n13948), .B1(n13947), .B2(n13946), .ZN(
        n13960) );
  NAND2_X1 U15458 ( .A1(n13950), .A2(n13949), .ZN(n13951) );
  NAND3_X1 U15459 ( .A1(n13952), .A2(n13973), .A3(n13951), .ZN(n13957) );
  AOI22_X1 U15460 ( .A1(n13955), .A2(n13967), .B1(n13954), .B2(n13953), .ZN(
        n13956) );
  AND2_X1 U15461 ( .A1(n13957), .A2(n13956), .ZN(n14054) );
  NOR2_X1 U15462 ( .A1(n14054), .A2(n13958), .ZN(n13959) );
  AOI211_X1 U15463 ( .C1(n13981), .C2(n13961), .A(n13960), .B(n13959), .ZN(
        n13962) );
  OAI21_X1 U15464 ( .B1(n14058), .B2(n13963), .A(n13962), .ZN(P3_U3220) );
  XNOR2_X1 U15465 ( .A(n13964), .B(n13966), .ZN(n14135) );
  INV_X1 U15466 ( .A(n14135), .ZN(n14064) );
  XNOR2_X1 U15467 ( .A(n13965), .B(n13966), .ZN(n13974) );
  NAND2_X1 U15468 ( .A1(n13968), .A2(n13967), .ZN(n13969) );
  OAI21_X1 U15469 ( .B1(n13971), .B2(n13970), .A(n13969), .ZN(n13972) );
  AOI21_X1 U15470 ( .B1(n13974), .B2(n13973), .A(n13972), .ZN(n13976) );
  NAND2_X1 U15471 ( .A1(n14135), .A2(n14052), .ZN(n13975) );
  MUX2_X1 U15472 ( .A(n13978), .B(n14132), .S(n13977), .Z(n13983) );
  AOI22_X1 U15473 ( .A1(n13981), .A2(n14060), .B1(n13980), .B2(n13979), .ZN(
        n13982) );
  OAI211_X1 U15474 ( .C1(n14064), .C2(n13984), .A(n13983), .B(n13982), .ZN(
        P3_U3221) );
  NAND2_X1 U15475 ( .A1(n16585), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13985) );
  NAND2_X1 U15476 ( .A1(n14065), .A2(n16587), .ZN(n13987) );
  OAI211_X1 U15477 ( .C1(n14067), .C2(n14051), .A(n13985), .B(n13987), .ZN(
        P3_U3490) );
  NAND2_X1 U15478 ( .A1(n16585), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n13986) );
  OAI211_X1 U15479 ( .C1(n14070), .C2(n14051), .A(n13987), .B(n13986), .ZN(
        P3_U3489) );
  NAND2_X1 U15480 ( .A1(n13988), .A2(n16578), .ZN(n13989) );
  NAND2_X1 U15481 ( .A1(n13990), .A2(n13989), .ZN(n14071) );
  INV_X1 U15482 ( .A(n13991), .ZN(n13992) );
  OAI21_X1 U15483 ( .B1(n14074), .B2(n14051), .A(n13992), .ZN(P3_U3487) );
  MUX2_X1 U15484 ( .A(n14075), .B(P3_REG1_REG_27__SCAN_IN), .S(n16585), .Z(
        n13994) );
  OAI22_X1 U15485 ( .A1(n13747), .A2(n14063), .B1(n14076), .B2(n14051), .ZN(
        n13993) );
  INV_X1 U15486 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13995) );
  MUX2_X1 U15487 ( .A(n13995), .B(n14079), .S(n16587), .Z(n13998) );
  NAND2_X1 U15488 ( .A1(n13996), .A2(n10089), .ZN(n13997) );
  OAI211_X1 U15489 ( .C1(n13999), .C2(n14063), .A(n13998), .B(n13997), .ZN(
        P3_U3485) );
  INV_X1 U15490 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n14002) );
  AOI21_X1 U15491 ( .B1(n14040), .B2(n14001), .A(n14000), .ZN(n14086) );
  MUX2_X1 U15492 ( .A(n14002), .B(n14086), .S(n16587), .Z(n14003) );
  OAI21_X1 U15493 ( .B1(n14089), .B2(n14063), .A(n14003), .ZN(P3_U3484) );
  MUX2_X1 U15494 ( .A(n14090), .B(P3_REG1_REG_24__SCAN_IN), .S(n16585), .Z(
        n14005) );
  OAI22_X1 U15495 ( .A1(n14092), .A2(n14063), .B1(n14091), .B2(n14051), .ZN(
        n14004) );
  OR2_X1 U15496 ( .A1(n14005), .A2(n14004), .ZN(P3_U3483) );
  INV_X1 U15497 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n14010) );
  INV_X1 U15498 ( .A(n16578), .ZN(n14034) );
  NOR2_X1 U15499 ( .A1(n14006), .A2(n14034), .ZN(n14009) );
  AOI21_X1 U15500 ( .B1(n14009), .B2(n14008), .A(n14007), .ZN(n14095) );
  MUX2_X1 U15501 ( .A(n14010), .B(n14095), .S(n16587), .Z(n14011) );
  OAI21_X1 U15502 ( .B1(n14098), .B2(n14051), .A(n14011), .ZN(P3_U3482) );
  NAND2_X1 U15503 ( .A1(n14012), .A2(n14040), .ZN(n14013) );
  OAI211_X1 U15504 ( .C1(n14015), .C2(n14102), .A(n14014), .B(n14013), .ZN(
        n14099) );
  MUX2_X1 U15505 ( .A(P3_REG1_REG_22__SCAN_IN), .B(n14099), .S(n16587), .Z(
        n14016) );
  INV_X1 U15506 ( .A(n14016), .ZN(n14017) );
  OAI21_X1 U15507 ( .B1(n14102), .B2(n14063), .A(n14017), .ZN(P3_U3481) );
  INV_X1 U15508 ( .A(n14018), .ZN(n14106) );
  INV_X1 U15509 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n14021) );
  AOI21_X1 U15510 ( .B1(n14040), .B2(n14020), .A(n14019), .ZN(n14103) );
  MUX2_X1 U15511 ( .A(n14021), .B(n14103), .S(n16587), .Z(n14022) );
  OAI21_X1 U15512 ( .B1(n14106), .B2(n14063), .A(n14022), .ZN(P3_U3480) );
  MUX2_X1 U15513 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n14107), .S(n16587), .Z(
        n14025) );
  INV_X1 U15514 ( .A(n14023), .ZN(n14108) );
  OAI22_X1 U15515 ( .A1(n14110), .A2(n14063), .B1(n14108), .B2(n14051), .ZN(
        n14024) );
  OR2_X1 U15516 ( .A1(n14025), .A2(n14024), .ZN(P3_U3479) );
  AOI21_X1 U15517 ( .B1(n14040), .B2(n14027), .A(n14026), .ZN(n14028) );
  OAI21_X1 U15518 ( .B1(n14034), .B2(n14029), .A(n14028), .ZN(n14113) );
  MUX2_X1 U15519 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n14113), .S(n16587), .Z(
        P3_U3478) );
  AOI21_X1 U15520 ( .B1(n14040), .B2(n14031), .A(n14030), .ZN(n14032) );
  OAI21_X1 U15521 ( .B1(n14034), .B2(n14033), .A(n14032), .ZN(n14114) );
  MUX2_X1 U15522 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n14114), .S(n16587), .Z(
        P3_U3477) );
  AOI21_X1 U15523 ( .B1(n14036), .B2(n16578), .A(n14035), .ZN(n14115) );
  MUX2_X1 U15524 ( .A(n14037), .B(n14115), .S(n16587), .Z(n14038) );
  OAI21_X1 U15525 ( .B1(n14118), .B2(n14051), .A(n14038), .ZN(P3_U3476) );
  AOI22_X1 U15526 ( .A1(n14041), .A2(n16578), .B1(n14040), .B2(n14039), .ZN(
        n14042) );
  NAND2_X1 U15527 ( .A1(n14043), .A2(n14042), .ZN(n14119) );
  MUX2_X1 U15528 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n14119), .S(n16587), .Z(
        P3_U3475) );
  AOI21_X1 U15529 ( .B1(n14045), .B2(n16578), .A(n14044), .ZN(n14120) );
  MUX2_X1 U15530 ( .A(n16373), .B(n14120), .S(n16587), .Z(n14046) );
  OAI21_X1 U15531 ( .B1(n14123), .B2(n14051), .A(n14046), .ZN(P3_U3474) );
  AOI21_X1 U15532 ( .B1(n14048), .B2(n16578), .A(n14047), .ZN(n14124) );
  MUX2_X1 U15533 ( .A(n14049), .B(n14124), .S(n16587), .Z(n14050) );
  OAI21_X1 U15534 ( .B1(n14051), .B2(n14127), .A(n14050), .ZN(P3_U3473) );
  NAND2_X1 U15535 ( .A1(n14130), .A2(n14052), .ZN(n14053) );
  OAI211_X1 U15536 ( .C1(n16580), .C2(n14055), .A(n14054), .B(n14053), .ZN(
        n14128) );
  MUX2_X1 U15537 ( .A(P3_REG1_REG_13__SCAN_IN), .B(n14128), .S(n16587), .Z(
        n14056) );
  INV_X1 U15538 ( .A(n14056), .ZN(n14057) );
  OAI21_X1 U15539 ( .B1(n14058), .B2(n14063), .A(n14057), .ZN(P3_U3472) );
  INV_X1 U15540 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14059) );
  MUX2_X1 U15541 ( .A(n14059), .B(n14132), .S(n16587), .Z(n14062) );
  NAND2_X1 U15542 ( .A1(n10089), .A2(n14060), .ZN(n14061) );
  OAI211_X1 U15543 ( .C1(n14064), .C2(n14063), .A(n14062), .B(n14061), .ZN(
        P3_U3471) );
  NAND2_X1 U15544 ( .A1(n16588), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n14066) );
  NAND2_X1 U15545 ( .A1(n14065), .A2(n16590), .ZN(n14069) );
  OAI211_X1 U15546 ( .C1(n14067), .C2(n14139), .A(n14066), .B(n14069), .ZN(
        P3_U3458) );
  NAND2_X1 U15547 ( .A1(n16588), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n14068) );
  OAI211_X1 U15548 ( .C1(n14070), .C2(n14139), .A(n14069), .B(n14068), .ZN(
        P3_U3457) );
  INV_X1 U15549 ( .A(n14072), .ZN(n14073) );
  OAI21_X1 U15550 ( .B1(n14074), .B2(n14139), .A(n14073), .ZN(P3_U3455) );
  MUX2_X1 U15551 ( .A(n14075), .B(P3_REG0_REG_27__SCAN_IN), .S(n16588), .Z(
        n14078) );
  OAI22_X1 U15552 ( .A1(n13747), .A2(n14109), .B1(n14076), .B2(n14139), .ZN(
        n14077) );
  INV_X1 U15553 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n14080) );
  MUX2_X1 U15554 ( .A(n14080), .B(n14079), .S(n16590), .Z(n14085) );
  NOR2_X1 U15555 ( .A1(n14081), .A2(n14139), .ZN(n14082) );
  AOI21_X1 U15556 ( .B1(n14083), .B2(n14134), .A(n14082), .ZN(n14084) );
  NAND2_X1 U15557 ( .A1(n14085), .A2(n14084), .ZN(P3_U3453) );
  INV_X1 U15558 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n14087) );
  MUX2_X1 U15559 ( .A(n14087), .B(n14086), .S(n16590), .Z(n14088) );
  OAI21_X1 U15560 ( .B1(n14089), .B2(n14109), .A(n14088), .ZN(P3_U3452) );
  MUX2_X1 U15561 ( .A(n14090), .B(P3_REG0_REG_24__SCAN_IN), .S(n16588), .Z(
        n14094) );
  OAI22_X1 U15562 ( .A1(n14092), .A2(n14109), .B1(n14091), .B2(n14139), .ZN(
        n14093) );
  OR2_X1 U15563 ( .A1(n14094), .A2(n14093), .ZN(P3_U3451) );
  INV_X1 U15564 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n14096) );
  MUX2_X1 U15565 ( .A(n14096), .B(n14095), .S(n16590), .Z(n14097) );
  OAI21_X1 U15566 ( .B1(n14098), .B2(n14139), .A(n14097), .ZN(P3_U3450) );
  MUX2_X1 U15567 ( .A(P3_REG0_REG_22__SCAN_IN), .B(n14099), .S(n16590), .Z(
        n14100) );
  INV_X1 U15568 ( .A(n14100), .ZN(n14101) );
  OAI21_X1 U15569 ( .B1(n14102), .B2(n14109), .A(n14101), .ZN(P3_U3449) );
  INV_X1 U15570 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n14104) );
  MUX2_X1 U15571 ( .A(n14104), .B(n14103), .S(n16590), .Z(n14105) );
  OAI21_X1 U15572 ( .B1(n14106), .B2(n14109), .A(n14105), .ZN(P3_U3448) );
  MUX2_X1 U15573 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n14107), .S(n16590), .Z(
        n14112) );
  OAI22_X1 U15574 ( .A1(n14110), .A2(n14109), .B1(n14108), .B2(n14139), .ZN(
        n14111) );
  OR2_X1 U15575 ( .A1(n14112), .A2(n14111), .ZN(P3_U3447) );
  MUX2_X1 U15576 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n14113), .S(n16590), .Z(
        P3_U3446) );
  MUX2_X1 U15577 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n14114), .S(n16590), .Z(
        P3_U3444) );
  MUX2_X1 U15578 ( .A(n14116), .B(n14115), .S(n16590), .Z(n14117) );
  OAI21_X1 U15579 ( .B1(n14118), .B2(n14139), .A(n14117), .ZN(P3_U3441) );
  MUX2_X1 U15580 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n14119), .S(n16590), .Z(
        P3_U3438) );
  INV_X1 U15581 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n14121) );
  MUX2_X1 U15582 ( .A(n14121), .B(n14120), .S(n16590), .Z(n14122) );
  OAI21_X1 U15583 ( .B1(n14123), .B2(n14139), .A(n14122), .ZN(P3_U3435) );
  MUX2_X1 U15584 ( .A(n14125), .B(n14124), .S(n16590), .Z(n14126) );
  OAI21_X1 U15585 ( .B1(n14139), .B2(n14127), .A(n14126), .ZN(P3_U3432) );
  MUX2_X1 U15586 ( .A(P3_REG0_REG_13__SCAN_IN), .B(n14128), .S(n16590), .Z(
        n14129) );
  AOI21_X1 U15587 ( .B1(n14134), .B2(n14130), .A(n14129), .ZN(n14131) );
  INV_X1 U15588 ( .A(n14131), .ZN(P3_U3429) );
  INV_X1 U15589 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14133) );
  MUX2_X1 U15590 ( .A(n14133), .B(n14132), .S(n16590), .Z(n14137) );
  NAND2_X1 U15591 ( .A1(n14135), .A2(n14134), .ZN(n14136) );
  OAI211_X1 U15592 ( .C1(n14139), .C2(n14138), .A(n14137), .B(n14136), .ZN(
        P3_U3426) );
  MUX2_X1 U15593 ( .A(P3_D_REG_1__SCAN_IN), .B(n14141), .S(n14140), .Z(
        P3_U3377) );
  INV_X1 U15594 ( .A(n14142), .ZN(n14148) );
  NOR4_X1 U15595 ( .A1(n14144), .A2(P3_IR_REG_30__SCAN_IN), .A3(n14143), .A4(
        P3_U3151), .ZN(n14145) );
  AOI21_X1 U15596 ( .B1(SI_31_), .B2(n14146), .A(n14145), .ZN(n14147) );
  OAI21_X1 U15597 ( .B1(n14148), .B2(n14154), .A(n14147), .ZN(P3_U3264) );
  INV_X1 U15598 ( .A(n14149), .ZN(n14153) );
  INV_X1 U15599 ( .A(SI_29_), .ZN(n14151) );
  MUX2_X1 U15600 ( .A(n14156), .B(n14155), .S(P3_STATE_REG_SCAN_IN), .Z(
        P3_U3294) );
  NAND2_X1 U15601 ( .A1(n14671), .A2(n14914), .ZN(n14160) );
  NAND2_X1 U15602 ( .A1(n14157), .A2(n14707), .ZN(n14159) );
  MUX2_X1 U15603 ( .A(n14160), .B(n14159), .S(n14158), .Z(n14165) );
  OAI22_X1 U15604 ( .A1(n14870), .A2(n14953), .B1(n14942), .B2(n14951), .ZN(
        n14897) );
  INV_X1 U15605 ( .A(n14897), .ZN(n14162) );
  OAI22_X1 U15606 ( .A1(n14162), .A2(n14650), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14161), .ZN(n14163) );
  AOI21_X1 U15607 ( .B1(n14904), .B2(n14700), .A(n14163), .ZN(n14164) );
  OAI211_X1 U15608 ( .C1(n7952), .C2(n14705), .A(n14165), .B(n14164), .ZN(
        P2_U3188) );
  AOI21_X1 U15609 ( .B1(n14167), .B2(n14166), .A(n14686), .ZN(n14169) );
  NAND2_X1 U15610 ( .A1(n14169), .A2(n14168), .ZN(n14174) );
  AOI22_X1 U15611 ( .A1(n14681), .A2(n14171), .B1(n14691), .B2(n14170), .ZN(
        n14173) );
  MUX2_X1 U15612 ( .A(n14683), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n14172) );
  NAND3_X1 U15613 ( .A1(n14174), .A2(n14173), .A3(n14172), .ZN(P2_U3190) );
  INV_X1 U15614 ( .A(n15057), .ZN(n14975) );
  INV_X1 U15615 ( .A(n14175), .ZN(n14176) );
  AOI21_X1 U15616 ( .B1(n14176), .B2(n14684), .A(n14686), .ZN(n14180) );
  NOR3_X1 U15617 ( .A1(n14178), .A2(n14177), .A3(n14694), .ZN(n14179) );
  OAI21_X1 U15618 ( .B1(n14180), .B2(n14179), .A(n14660), .ZN(n14186) );
  NAND2_X1 U15619 ( .A1(n14716), .A2(n14913), .ZN(n14182) );
  NAND2_X1 U15620 ( .A1(n14718), .A2(n14911), .ZN(n14181) );
  NAND2_X1 U15621 ( .A1(n14182), .A2(n14181), .ZN(n14965) );
  NOR2_X1 U15622 ( .A1(n14683), .A2(n14971), .ZN(n14183) );
  AOI211_X1 U15623 ( .C1(n14681), .C2(n14965), .A(n14184), .B(n14183), .ZN(
        n14185) );
  OAI211_X1 U15624 ( .C1(n14975), .C2(n14705), .A(n14186), .B(n14185), .ZN(
        P2_U3191) );
  INV_X1 U15625 ( .A(n14861), .ZN(n14819) );
  NOR3_X1 U15626 ( .A1(n14187), .A2(n14819), .A3(n14694), .ZN(n14188) );
  AOI21_X1 U15627 ( .B1(n14189), .B2(n14707), .A(n14188), .ZN(n14200) );
  INV_X1 U15628 ( .A(n15011), .ZN(n14827) );
  MUX2_X1 U15629 ( .A(n14822), .B(n14827), .S(n14930), .Z(n14191) );
  XNOR2_X1 U15630 ( .A(n14191), .B(n14190), .ZN(n14199) );
  INV_X1 U15631 ( .A(n14194), .ZN(n14825) );
  AOI22_X1 U15632 ( .A1(n14825), .A2(n14700), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14197) );
  AOI22_X1 U15633 ( .A1(n14713), .A2(n14702), .B1(n14861), .B2(n14701), .ZN(
        n14196) );
  NAND2_X1 U15634 ( .A1(n15011), .A2(n14691), .ZN(n14195) );
  OAI21_X1 U15635 ( .B1(n14200), .B2(n14199), .A(n14198), .ZN(P2_U3192) );
  AOI22_X1 U15636 ( .A1(n14671), .A2(n14202), .B1(n14707), .B2(n14201), .ZN(
        n14209) );
  AOI22_X1 U15637 ( .A1(n14681), .A2(n14204), .B1(n14707), .B2(n14203), .ZN(
        n14207) );
  AOI22_X1 U15638 ( .A1(n16420), .A2(n14691), .B1(n14205), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n14206) );
  OAI211_X1 U15639 ( .C1(n14209), .C2(n14208), .A(n14207), .B(n14206), .ZN(
        n14615) );
  XOR2_X1 U15640 ( .A(SI_30_), .B(keyinput_130), .Z(n14212) );
  XNOR2_X1 U15641 ( .A(n14407), .B(keyinput_132), .ZN(n14211) );
  XNOR2_X1 U15642 ( .A(SI_31_), .B(keyinput_129), .ZN(n14210) );
  NOR3_X1 U15643 ( .A1(n14212), .A2(n14211), .A3(n14210), .ZN(n14215) );
  XOR2_X1 U15644 ( .A(SI_29_), .B(keyinput_131), .Z(n14214) );
  XOR2_X1 U15645 ( .A(keyinput_128), .B(P3_WR_REG_SCAN_IN), .Z(n14213) );
  NAND3_X1 U15646 ( .A1(n14215), .A2(n14214), .A3(n14213), .ZN(n14218) );
  XOR2_X1 U15647 ( .A(SI_27_), .B(keyinput_133), .Z(n14217) );
  XNOR2_X1 U15648 ( .A(SI_26_), .B(keyinput_134), .ZN(n14216) );
  AOI21_X1 U15649 ( .B1(n14218), .B2(n14217), .A(n14216), .ZN(n14221) );
  XNOR2_X1 U15650 ( .A(SI_24_), .B(keyinput_136), .ZN(n14220) );
  XNOR2_X1 U15651 ( .A(SI_25_), .B(keyinput_135), .ZN(n14219) );
  NOR3_X1 U15652 ( .A1(n14221), .A2(n14220), .A3(n14219), .ZN(n14224) );
  XOR2_X1 U15653 ( .A(SI_23_), .B(keyinput_137), .Z(n14223) );
  XNOR2_X1 U15654 ( .A(n14417), .B(keyinput_138), .ZN(n14222) );
  OAI21_X1 U15655 ( .B1(n14224), .B2(n14223), .A(n14222), .ZN(n14227) );
  XOR2_X1 U15656 ( .A(SI_21_), .B(keyinput_139), .Z(n14226) );
  XNOR2_X1 U15657 ( .A(SI_20_), .B(keyinput_140), .ZN(n14225) );
  NAND3_X1 U15658 ( .A1(n14227), .A2(n14226), .A3(n14225), .ZN(n14230) );
  XNOR2_X1 U15659 ( .A(n14425), .B(keyinput_142), .ZN(n14229) );
  XNOR2_X1 U15660 ( .A(SI_19_), .B(keyinput_141), .ZN(n14228) );
  NAND3_X1 U15661 ( .A1(n14230), .A2(n14229), .A3(n14228), .ZN(n14234) );
  XNOR2_X1 U15662 ( .A(n14430), .B(keyinput_145), .ZN(n14233) );
  XNOR2_X1 U15663 ( .A(SI_17_), .B(keyinput_143), .ZN(n14232) );
  XNOR2_X1 U15664 ( .A(SI_16_), .B(keyinput_144), .ZN(n14231) );
  NAND4_X1 U15665 ( .A1(n14234), .A2(n14233), .A3(n14232), .A4(n14231), .ZN(
        n14242) );
  XNOR2_X1 U15666 ( .A(n14235), .B(keyinput_149), .ZN(n14240) );
  XNOR2_X1 U15667 ( .A(n14236), .B(keyinput_148), .ZN(n14239) );
  XNOR2_X1 U15668 ( .A(n14435), .B(keyinput_146), .ZN(n14238) );
  XNOR2_X1 U15669 ( .A(SI_13_), .B(keyinput_147), .ZN(n14237) );
  NOR4_X1 U15670 ( .A1(n14240), .A2(n14239), .A3(n14238), .A4(n14237), .ZN(
        n14241) );
  NAND2_X1 U15671 ( .A1(n14242), .A2(n14241), .ZN(n14246) );
  XOR2_X1 U15672 ( .A(SI_8_), .B(keyinput_152), .Z(n14245) );
  XNOR2_X1 U15673 ( .A(n14440), .B(keyinput_150), .ZN(n14244) );
  XNOR2_X1 U15674 ( .A(SI_9_), .B(keyinput_151), .ZN(n14243) );
  NAND4_X1 U15675 ( .A1(n14246), .A2(n14245), .A3(n14244), .A4(n14243), .ZN(
        n14250) );
  XNOR2_X1 U15676 ( .A(SI_7_), .B(keyinput_153), .ZN(n14249) );
  XOR2_X1 U15677 ( .A(SI_6_), .B(keyinput_154), .Z(n14248) );
  XNOR2_X1 U15678 ( .A(SI_5_), .B(keyinput_155), .ZN(n14247) );
  AOI211_X1 U15679 ( .C1(n14250), .C2(n14249), .A(n14248), .B(n14247), .ZN(
        n14253) );
  XNOR2_X1 U15680 ( .A(SI_4_), .B(keyinput_156), .ZN(n14252) );
  XNOR2_X1 U15681 ( .A(SI_3_), .B(keyinput_157), .ZN(n14251) );
  NOR3_X1 U15682 ( .A1(n14253), .A2(n14252), .A3(n14251), .ZN(n14256) );
  XOR2_X1 U15683 ( .A(SI_2_), .B(keyinput_158), .Z(n14255) );
  XOR2_X1 U15684 ( .A(SI_1_), .B(keyinput_159), .Z(n14254) );
  NOR3_X1 U15685 ( .A1(n14256), .A2(n14255), .A3(n14254), .ZN(n14260) );
  XNOR2_X1 U15686 ( .A(SI_0_), .B(keyinput_160), .ZN(n14259) );
  INV_X1 U15687 ( .A(P3_RD_REG_SCAN_IN), .ZN(n16384) );
  XNOR2_X1 U15688 ( .A(n16384), .B(keyinput_161), .ZN(n14258) );
  XNOR2_X1 U15689 ( .A(P3_U3151), .B(keyinput_162), .ZN(n14257) );
  OAI211_X1 U15690 ( .C1(n14260), .C2(n14259), .A(n14258), .B(n14257), .ZN(
        n14263) );
  XOR2_X1 U15691 ( .A(P3_REG3_REG_7__SCAN_IN), .B(keyinput_163), .Z(n14262) );
  XNOR2_X1 U15692 ( .A(P3_REG3_REG_27__SCAN_IN), .B(keyinput_164), .ZN(n14261)
         );
  AOI21_X1 U15693 ( .B1(n14263), .B2(n14262), .A(n14261), .ZN(n14266) );
  XNOR2_X1 U15694 ( .A(n14464), .B(keyinput_165), .ZN(n14265) );
  XOR2_X1 U15695 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput_166), .Z(n14264)
         );
  OAI21_X1 U15696 ( .B1(n14266), .B2(n14265), .A(n14264), .ZN(n14280) );
  AOI22_X1 U15697 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_172), .B1(
        P3_REG3_REG_19__SCAN_IN), .B2(keyinput_169), .ZN(n14267) );
  OAI221_X1 U15698 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_172), .C1(
        P3_REG3_REG_19__SCAN_IN), .C2(keyinput_169), .A(n14267), .ZN(n14270)
         );
  XNOR2_X1 U15699 ( .A(P3_REG3_REG_25__SCAN_IN), .B(keyinput_175), .ZN(n14269)
         );
  XNOR2_X1 U15700 ( .A(P3_REG3_REG_21__SCAN_IN), .B(keyinput_173), .ZN(n14268)
         );
  NOR3_X1 U15701 ( .A1(n14270), .A2(n14269), .A3(n14268), .ZN(n14279) );
  AOI22_X1 U15702 ( .A1(P3_REG3_REG_28__SCAN_IN), .A2(keyinput_170), .B1(
        n14272), .B2(keyinput_167), .ZN(n14271) );
  OAI221_X1 U15703 ( .B1(P3_REG3_REG_28__SCAN_IN), .B2(keyinput_170), .C1(
        n14272), .C2(keyinput_167), .A(n14271), .ZN(n14277) );
  XNOR2_X1 U15704 ( .A(n14273), .B(keyinput_171), .ZN(n14276) );
  XNOR2_X1 U15705 ( .A(n14472), .B(keyinput_168), .ZN(n14275) );
  XNOR2_X1 U15706 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput_174), .ZN(n14274)
         );
  NOR4_X1 U15707 ( .A1(n14277), .A2(n14276), .A3(n14275), .A4(n14274), .ZN(
        n14278) );
  NAND3_X1 U15708 ( .A1(n14280), .A2(n14279), .A3(n14278), .ZN(n14287) );
  XOR2_X1 U15709 ( .A(P3_REG3_REG_17__SCAN_IN), .B(keyinput_178), .Z(n14283)
         );
  XNOR2_X1 U15710 ( .A(P3_REG3_REG_5__SCAN_IN), .B(keyinput_177), .ZN(n14282)
         );
  XNOR2_X1 U15711 ( .A(P3_REG3_REG_16__SCAN_IN), .B(keyinput_176), .ZN(n14281)
         );
  NOR3_X1 U15712 ( .A1(n14283), .A2(n14282), .A3(n14281), .ZN(n14286) );
  XOR2_X1 U15713 ( .A(P3_REG3_REG_24__SCAN_IN), .B(keyinput_179), .Z(n14285)
         );
  XNOR2_X1 U15714 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput_180), .ZN(n14284)
         );
  AOI211_X1 U15715 ( .C1(n14287), .C2(n14286), .A(n14285), .B(n14284), .ZN(
        n14290) );
  XNOR2_X1 U15716 ( .A(P3_REG3_REG_9__SCAN_IN), .B(keyinput_181), .ZN(n14289)
         );
  XNOR2_X1 U15717 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_182), .ZN(n14288)
         );
  OAI21_X1 U15718 ( .B1(n14290), .B2(n14289), .A(n14288), .ZN(n14294) );
  XNOR2_X1 U15719 ( .A(n14291), .B(keyinput_183), .ZN(n14293) );
  XNOR2_X1 U15720 ( .A(P3_REG3_REG_13__SCAN_IN), .B(keyinput_184), .ZN(n14292)
         );
  NAND3_X1 U15721 ( .A1(n14294), .A2(n14293), .A3(n14292), .ZN(n14302) );
  XOR2_X1 U15722 ( .A(P3_REG3_REG_2__SCAN_IN), .B(keyinput_187), .Z(n14299) );
  XOR2_X1 U15723 ( .A(P3_REG3_REG_11__SCAN_IN), .B(keyinput_186), .Z(n14298)
         );
  XNOR2_X1 U15724 ( .A(n14295), .B(keyinput_188), .ZN(n14297) );
  XNOR2_X1 U15725 ( .A(P3_REG3_REG_22__SCAN_IN), .B(keyinput_185), .ZN(n14296)
         );
  NOR4_X1 U15726 ( .A1(n14299), .A2(n14298), .A3(n14297), .A4(n14296), .ZN(
        n14301) );
  XOR2_X1 U15727 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput_189), .Z(n14300) );
  AOI21_X1 U15728 ( .B1(n14302), .B2(n14301), .A(n14300), .ZN(n14305) );
  XNOR2_X1 U15729 ( .A(n14505), .B(keyinput_190), .ZN(n14304) );
  XOR2_X1 U15730 ( .A(P3_REG3_REG_15__SCAN_IN), .B(keyinput_191), .Z(n14303)
         );
  OAI21_X1 U15731 ( .B1(n14305), .B2(n14304), .A(n14303), .ZN(n14311) );
  XOR2_X1 U15732 ( .A(P3_B_REG_SCAN_IN), .B(keyinput_192), .Z(n14310) );
  XOR2_X1 U15733 ( .A(keyinput_195), .B(P3_DATAO_REG_29__SCAN_IN), .Z(n14308)
         );
  XOR2_X1 U15734 ( .A(keyinput_194), .B(P3_DATAO_REG_30__SCAN_IN), .Z(n14307)
         );
  XNOR2_X1 U15735 ( .A(keyinput_193), .B(P3_DATAO_REG_31__SCAN_IN), .ZN(n14306) );
  NAND3_X1 U15736 ( .A1(n14308), .A2(n14307), .A3(n14306), .ZN(n14309) );
  AOI21_X1 U15737 ( .B1(n14311), .B2(n14310), .A(n14309), .ZN(n14314) );
  XNOR2_X1 U15738 ( .A(keyinput_197), .B(P3_DATAO_REG_27__SCAN_IN), .ZN(n14313) );
  XNOR2_X1 U15739 ( .A(keyinput_196), .B(P3_DATAO_REG_28__SCAN_IN), .ZN(n14312) );
  NOR3_X1 U15740 ( .A1(n14314), .A2(n14313), .A3(n14312), .ZN(n14317) );
  XNOR2_X1 U15741 ( .A(keyinput_198), .B(P3_DATAO_REG_26__SCAN_IN), .ZN(n14316) );
  XOR2_X1 U15742 ( .A(keyinput_199), .B(P3_DATAO_REG_25__SCAN_IN), .Z(n14315)
         );
  OAI21_X1 U15743 ( .B1(n14317), .B2(n14316), .A(n14315), .ZN(n14320) );
  XOR2_X1 U15744 ( .A(keyinput_201), .B(P3_DATAO_REG_23__SCAN_IN), .Z(n14319)
         );
  XNOR2_X1 U15745 ( .A(keyinput_200), .B(P3_DATAO_REG_24__SCAN_IN), .ZN(n14318) );
  NAND3_X1 U15746 ( .A1(n14320), .A2(n14319), .A3(n14318), .ZN(n14324) );
  XNOR2_X1 U15747 ( .A(keyinput_202), .B(P3_DATAO_REG_22__SCAN_IN), .ZN(n14323) );
  XOR2_X1 U15748 ( .A(keyinput_203), .B(P3_DATAO_REG_21__SCAN_IN), .Z(n14322)
         );
  XNOR2_X1 U15749 ( .A(keyinput_204), .B(P3_DATAO_REG_20__SCAN_IN), .ZN(n14321) );
  AOI211_X1 U15750 ( .C1(n14324), .C2(n14323), .A(n14322), .B(n14321), .ZN(
        n14327) );
  XOR2_X1 U15751 ( .A(keyinput_205), .B(P3_DATAO_REG_19__SCAN_IN), .Z(n14326)
         );
  XOR2_X1 U15752 ( .A(keyinput_206), .B(P3_DATAO_REG_18__SCAN_IN), .Z(n14325)
         );
  NOR3_X1 U15753 ( .A1(n14327), .A2(n14326), .A3(n14325), .ZN(n14343) );
  INV_X1 U15754 ( .A(keyinput_208), .ZN(n14334) );
  INV_X1 U15755 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n14534) );
  INV_X1 U15756 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n14328) );
  OAI22_X1 U15757 ( .A1(n14534), .A2(keyinput_210), .B1(n14328), .B2(
        keyinput_208), .ZN(n14331) );
  INV_X1 U15758 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n14533) );
  OAI22_X1 U15759 ( .A1(n14533), .A2(keyinput_209), .B1(
        P3_DATAO_REG_11__SCAN_IN), .B2(keyinput_213), .ZN(n14330) );
  INV_X1 U15760 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n14336) );
  OAI22_X1 U15761 ( .A1(n14336), .A2(keyinput_212), .B1(
        P3_DATAO_REG_13__SCAN_IN), .B2(keyinput_211), .ZN(n14329) );
  NOR3_X1 U15762 ( .A1(n14331), .A2(n14330), .A3(n14329), .ZN(n14333) );
  NAND2_X1 U15763 ( .A1(P3_DATAO_REG_11__SCAN_IN), .A2(keyinput_213), .ZN(
        n14332) );
  OAI211_X1 U15764 ( .C1(n14334), .C2(P3_DATAO_REG_16__SCAN_IN), .A(n14333), 
        .B(n14332), .ZN(n14335) );
  INV_X1 U15765 ( .A(n14335), .ZN(n14340) );
  AOI22_X1 U15766 ( .A1(keyinput_212), .A2(n14336), .B1(n14534), .B2(
        keyinput_210), .ZN(n14339) );
  AOI22_X1 U15767 ( .A1(n14533), .A2(keyinput_209), .B1(keyinput_211), .B2(
        P3_DATAO_REG_13__SCAN_IN), .ZN(n14338) );
  XNOR2_X1 U15768 ( .A(keyinput_207), .B(P3_DATAO_REG_17__SCAN_IN), .ZN(n14337) );
  NAND4_X1 U15769 ( .A1(n14340), .A2(n14339), .A3(n14338), .A4(n14337), .ZN(
        n14342) );
  XOR2_X1 U15770 ( .A(keyinput_214), .B(P3_DATAO_REG_10__SCAN_IN), .Z(n14341)
         );
  OAI21_X1 U15771 ( .B1(n14343), .B2(n14342), .A(n14341), .ZN(n14353) );
  XOR2_X1 U15772 ( .A(keyinput_218), .B(P3_DATAO_REG_6__SCAN_IN), .Z(n14347)
         );
  XOR2_X1 U15773 ( .A(keyinput_216), .B(P3_DATAO_REG_8__SCAN_IN), .Z(n14346)
         );
  XNOR2_X1 U15774 ( .A(keyinput_215), .B(P3_DATAO_REG_9__SCAN_IN), .ZN(n14345)
         );
  XNOR2_X1 U15775 ( .A(keyinput_217), .B(P3_DATAO_REG_7__SCAN_IN), .ZN(n14344)
         );
  NOR4_X1 U15776 ( .A1(n14347), .A2(n14346), .A3(n14345), .A4(n14344), .ZN(
        n14352) );
  XOR2_X1 U15777 ( .A(keyinput_220), .B(P3_DATAO_REG_4__SCAN_IN), .Z(n14350)
         );
  XOR2_X1 U15778 ( .A(keyinput_221), .B(P3_DATAO_REG_3__SCAN_IN), .Z(n14349)
         );
  XOR2_X1 U15779 ( .A(keyinput_219), .B(P3_DATAO_REG_5__SCAN_IN), .Z(n14348)
         );
  NAND3_X1 U15780 ( .A1(n14350), .A2(n14349), .A3(n14348), .ZN(n14351) );
  AOI21_X1 U15781 ( .B1(n14353), .B2(n14352), .A(n14351), .ZN(n14356) );
  XNOR2_X1 U15782 ( .A(keyinput_223), .B(P3_DATAO_REG_1__SCAN_IN), .ZN(n14355)
         );
  XNOR2_X1 U15783 ( .A(keyinput_222), .B(P3_DATAO_REG_2__SCAN_IN), .ZN(n14354)
         );
  NOR3_X1 U15784 ( .A1(n14356), .A2(n14355), .A3(n14354), .ZN(n14359) );
  XNOR2_X1 U15785 ( .A(keyinput_224), .B(P3_DATAO_REG_0__SCAN_IN), .ZN(n14358)
         );
  XOR2_X1 U15786 ( .A(keyinput_225), .B(P3_ADDR_REG_0__SCAN_IN), .Z(n14357) );
  OAI21_X1 U15787 ( .B1(n14359), .B2(n14358), .A(n14357), .ZN(n14363) );
  XNOR2_X1 U15788 ( .A(keyinput_226), .B(P3_ADDR_REG_1__SCAN_IN), .ZN(n14362)
         );
  XOR2_X1 U15789 ( .A(keyinput_228), .B(P3_ADDR_REG_3__SCAN_IN), .Z(n14361) );
  XNOR2_X1 U15790 ( .A(keyinput_227), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n14360)
         );
  AOI211_X1 U15791 ( .C1(n14363), .C2(n14362), .A(n14361), .B(n14360), .ZN(
        n14367) );
  XOR2_X1 U15792 ( .A(keyinput_229), .B(P3_ADDR_REG_4__SCAN_IN), .Z(n14366) );
  XOR2_X1 U15793 ( .A(keyinput_231), .B(P3_ADDR_REG_6__SCAN_IN), .Z(n14365) );
  XOR2_X1 U15794 ( .A(keyinput_230), .B(P3_ADDR_REG_5__SCAN_IN), .Z(n14364) );
  OAI211_X1 U15795 ( .C1(n14367), .C2(n14366), .A(n14365), .B(n14364), .ZN(
        n14370) );
  XOR2_X1 U15796 ( .A(keyinput_232), .B(P3_ADDR_REG_7__SCAN_IN), .Z(n14369) );
  XNOR2_X1 U15797 ( .A(keyinput_233), .B(P3_ADDR_REG_8__SCAN_IN), .ZN(n14368)
         );
  AOI21_X1 U15798 ( .B1(n14370), .B2(n14369), .A(n14368), .ZN(n14373) );
  XOR2_X1 U15799 ( .A(keyinput_234), .B(P3_ADDR_REG_9__SCAN_IN), .Z(n14372) );
  XNOR2_X1 U15800 ( .A(n16160), .B(keyinput_235), .ZN(n14371) );
  OAI21_X1 U15801 ( .B1(n14373), .B2(n14372), .A(n14371), .ZN(n14376) );
  XOR2_X1 U15802 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_236), .Z(n14375) );
  XNOR2_X1 U15803 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_237), .ZN(n14374) );
  AOI21_X1 U15804 ( .B1(n14376), .B2(n14375), .A(n14374), .ZN(n14379) );
  XOR2_X1 U15805 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_238), .Z(n14378) );
  XNOR2_X1 U15806 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_239), .ZN(n14377) );
  OAI21_X1 U15807 ( .B1(n14379), .B2(n14378), .A(n14377), .ZN(n14384) );
  XNOR2_X1 U15808 ( .A(n14587), .B(keyinput_241), .ZN(n14383) );
  XOR2_X1 U15809 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_242), .Z(n14382) );
  XNOR2_X1 U15810 ( .A(n14380), .B(keyinput_240), .ZN(n14381) );
  NAND4_X1 U15811 ( .A1(n14384), .A2(n14383), .A3(n14382), .A4(n14381), .ZN(
        n14387) );
  XNOR2_X1 U15812 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_243), .ZN(n14386) );
  XNOR2_X1 U15813 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_244), .ZN(n14385) );
  AOI21_X1 U15814 ( .B1(n14387), .B2(n14386), .A(n14385), .ZN(n14390) );
  XNOR2_X1 U15815 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_245), .ZN(n14389)
         );
  XNOR2_X1 U15816 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_246), .ZN(n14388)
         );
  OAI21_X1 U15817 ( .B1(n14390), .B2(n14389), .A(n14388), .ZN(n14396) );
  XNOR2_X1 U15818 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_248), .ZN(n14392)
         );
  XNOR2_X1 U15819 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_249), .ZN(n14391)
         );
  NOR2_X1 U15820 ( .A1(n14392), .A2(n14391), .ZN(n14395) );
  XNOR2_X1 U15821 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_250), .ZN(n14394)
         );
  XNOR2_X1 U15822 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_247), .ZN(n14393)
         );
  NAND4_X1 U15823 ( .A1(n14396), .A2(n14395), .A3(n14394), .A4(n14393), .ZN(
        n14403) );
  XOR2_X1 U15824 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_251), .Z(n14402) );
  XOR2_X1 U15825 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_254), .Z(n14400) );
  XNOR2_X1 U15826 ( .A(n14606), .B(keyinput_252), .ZN(n14399) );
  XNOR2_X1 U15827 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_255), .ZN(n14398)
         );
  XNOR2_X1 U15828 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_253), .ZN(n14397)
         );
  NAND4_X1 U15829 ( .A1(n14400), .A2(n14399), .A3(n14398), .A4(n14397), .ZN(
        n14401) );
  AOI21_X1 U15830 ( .B1(n14403), .B2(n14402), .A(n14401), .ZN(n14613) );
  XOR2_X1 U15831 ( .A(SI_31_), .B(keyinput_1), .Z(n14406) );
  XNOR2_X1 U15832 ( .A(SI_29_), .B(keyinput_3), .ZN(n14405) );
  XNOR2_X1 U15833 ( .A(SI_30_), .B(keyinput_2), .ZN(n14404) );
  NAND3_X1 U15834 ( .A1(n14406), .A2(n14405), .A3(n14404), .ZN(n14410) );
  XNOR2_X1 U15835 ( .A(n14407), .B(keyinput_4), .ZN(n14409) );
  XNOR2_X1 U15836 ( .A(P3_WR_REG_SCAN_IN), .B(keyinput_0), .ZN(n14408) );
  NOR3_X1 U15837 ( .A1(n14410), .A2(n14409), .A3(n14408), .ZN(n14413) );
  XOR2_X1 U15838 ( .A(SI_27_), .B(keyinput_5), .Z(n14412) );
  XOR2_X1 U15839 ( .A(SI_26_), .B(keyinput_6), .Z(n14411) );
  OAI21_X1 U15840 ( .B1(n14413), .B2(n14412), .A(n14411), .ZN(n14416) );
  XOR2_X1 U15841 ( .A(SI_24_), .B(keyinput_8), .Z(n14415) );
  XNOR2_X1 U15842 ( .A(SI_25_), .B(keyinput_7), .ZN(n14414) );
  NAND3_X1 U15843 ( .A1(n14416), .A2(n14415), .A3(n14414), .ZN(n14420) );
  XOR2_X1 U15844 ( .A(SI_23_), .B(keyinput_9), .Z(n14419) );
  XNOR2_X1 U15845 ( .A(n14417), .B(keyinput_10), .ZN(n14418) );
  AOI21_X1 U15846 ( .B1(n14420), .B2(n14419), .A(n14418), .ZN(n14423) );
  XOR2_X1 U15847 ( .A(SI_20_), .B(keyinput_12), .Z(n14422) );
  XOR2_X1 U15848 ( .A(SI_21_), .B(keyinput_11), .Z(n14421) );
  NOR3_X1 U15849 ( .A1(n14423), .A2(n14422), .A3(n14421), .ZN(n14428) );
  XNOR2_X1 U15850 ( .A(n14424), .B(keyinput_13), .ZN(n14427) );
  XNOR2_X1 U15851 ( .A(n14425), .B(keyinput_14), .ZN(n14426) );
  NOR3_X1 U15852 ( .A1(n14428), .A2(n14427), .A3(n14426), .ZN(n14434) );
  XNOR2_X1 U15853 ( .A(n14429), .B(keyinput_16), .ZN(n14433) );
  XNOR2_X1 U15854 ( .A(n14430), .B(keyinput_17), .ZN(n14432) );
  XNOR2_X1 U15855 ( .A(SI_17_), .B(keyinput_15), .ZN(n14431) );
  NOR4_X1 U15856 ( .A1(n14434), .A2(n14433), .A3(n14432), .A4(n14431), .ZN(
        n14446) );
  XOR2_X1 U15857 ( .A(SI_13_), .B(keyinput_19), .Z(n14439) );
  XNOR2_X1 U15858 ( .A(n14435), .B(keyinput_18), .ZN(n14438) );
  XNOR2_X1 U15859 ( .A(SI_11_), .B(keyinput_21), .ZN(n14437) );
  XNOR2_X1 U15860 ( .A(SI_12_), .B(keyinput_20), .ZN(n14436) );
  NAND4_X1 U15861 ( .A1(n14439), .A2(n14438), .A3(n14437), .A4(n14436), .ZN(
        n14445) );
  XOR2_X1 U15862 ( .A(SI_9_), .B(keyinput_23), .Z(n14443) );
  XNOR2_X1 U15863 ( .A(n14440), .B(keyinput_22), .ZN(n14442) );
  XNOR2_X1 U15864 ( .A(SI_8_), .B(keyinput_24), .ZN(n14441) );
  NOR3_X1 U15865 ( .A1(n14443), .A2(n14442), .A3(n14441), .ZN(n14444) );
  OAI21_X1 U15866 ( .B1(n14446), .B2(n14445), .A(n14444), .ZN(n14450) );
  XNOR2_X1 U15867 ( .A(SI_7_), .B(keyinput_25), .ZN(n14449) );
  XOR2_X1 U15868 ( .A(SI_6_), .B(keyinput_26), .Z(n14448) );
  XNOR2_X1 U15869 ( .A(SI_5_), .B(keyinput_27), .ZN(n14447) );
  AOI211_X1 U15870 ( .C1(n14450), .C2(n14449), .A(n14448), .B(n14447), .ZN(
        n14453) );
  XOR2_X1 U15871 ( .A(SI_4_), .B(keyinput_28), .Z(n14452) );
  XOR2_X1 U15872 ( .A(SI_3_), .B(keyinput_29), .Z(n14451) );
  NOR3_X1 U15873 ( .A1(n14453), .A2(n14452), .A3(n14451), .ZN(n14456) );
  XNOR2_X1 U15874 ( .A(SI_2_), .B(keyinput_30), .ZN(n14455) );
  XNOR2_X1 U15875 ( .A(SI_1_), .B(keyinput_31), .ZN(n14454) );
  NOR3_X1 U15876 ( .A1(n14456), .A2(n14455), .A3(n14454), .ZN(n14460) );
  XNOR2_X1 U15877 ( .A(SI_0_), .B(keyinput_32), .ZN(n14459) );
  XNOR2_X1 U15878 ( .A(P3_RD_REG_SCAN_IN), .B(keyinput_33), .ZN(n14458) );
  XNOR2_X1 U15879 ( .A(P3_STATE_REG_SCAN_IN), .B(keyinput_34), .ZN(n14457) );
  OAI211_X1 U15880 ( .C1(n14460), .C2(n14459), .A(n14458), .B(n14457), .ZN(
        n14463) );
  XNOR2_X1 U15881 ( .A(P3_REG3_REG_7__SCAN_IN), .B(keyinput_35), .ZN(n14462)
         );
  XOR2_X1 U15882 ( .A(P3_REG3_REG_27__SCAN_IN), .B(keyinput_36), .Z(n14461) );
  AOI21_X1 U15883 ( .B1(n14463), .B2(n14462), .A(n14461), .ZN(n14467) );
  XNOR2_X1 U15884 ( .A(n14464), .B(keyinput_37), .ZN(n14466) );
  XNOR2_X1 U15885 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput_38), .ZN(n14465)
         );
  OAI21_X1 U15886 ( .B1(n14467), .B2(n14466), .A(n14465), .ZN(n14482) );
  OAI22_X1 U15887 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput_46), .B1(
        keyinput_43), .B2(P3_REG3_REG_8__SCAN_IN), .ZN(n14468) );
  AOI221_X1 U15888 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_46), .C1(
        P3_REG3_REG_8__SCAN_IN), .C2(keyinput_43), .A(n14468), .ZN(n14481) );
  OAI22_X1 U15889 ( .A1(n14470), .A2(keyinput_41), .B1(P3_REG3_REG_25__SCAN_IN), .B2(keyinput_47), .ZN(n14469) );
  AOI221_X1 U15890 ( .B1(n14470), .B2(keyinput_41), .C1(keyinput_47), .C2(
        P3_REG3_REG_25__SCAN_IN), .A(n14469), .ZN(n14471) );
  INV_X1 U15891 ( .A(n14471), .ZN(n14479) );
  XNOR2_X1 U15892 ( .A(P3_REG3_REG_21__SCAN_IN), .B(keyinput_45), .ZN(n14478)
         );
  XNOR2_X1 U15893 ( .A(P3_REG3_REG_10__SCAN_IN), .B(keyinput_39), .ZN(n14477)
         );
  XNOR2_X1 U15894 ( .A(n14472), .B(keyinput_40), .ZN(n14475) );
  XNOR2_X1 U15895 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_44), .ZN(n14474)
         );
  XNOR2_X1 U15896 ( .A(P3_REG3_REG_28__SCAN_IN), .B(keyinput_42), .ZN(n14473)
         );
  NAND3_X1 U15897 ( .A1(n14475), .A2(n14474), .A3(n14473), .ZN(n14476) );
  NOR4_X1 U15898 ( .A1(n14479), .A2(n14478), .A3(n14477), .A4(n14476), .ZN(
        n14480) );
  NAND3_X1 U15899 ( .A1(n14482), .A2(n14481), .A3(n14480), .ZN(n14486) );
  XOR2_X1 U15900 ( .A(P3_REG3_REG_17__SCAN_IN), .B(keyinput_50), .Z(n14485) );
  XNOR2_X1 U15901 ( .A(P3_REG3_REG_16__SCAN_IN), .B(keyinput_48), .ZN(n14484)
         );
  XNOR2_X1 U15902 ( .A(P3_REG3_REG_5__SCAN_IN), .B(keyinput_49), .ZN(n14483)
         );
  NAND4_X1 U15903 ( .A1(n14486), .A2(n14485), .A3(n14484), .A4(n14483), .ZN(
        n14489) );
  XNOR2_X1 U15904 ( .A(P3_REG3_REG_24__SCAN_IN), .B(keyinput_51), .ZN(n14488)
         );
  XNOR2_X1 U15905 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput_52), .ZN(n14487)
         );
  NAND3_X1 U15906 ( .A1(n14489), .A2(n14488), .A3(n14487), .ZN(n14492) );
  XNOR2_X1 U15907 ( .A(P3_REG3_REG_9__SCAN_IN), .B(keyinput_53), .ZN(n14491)
         );
  XOR2_X1 U15908 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_54), .Z(n14490) );
  AOI21_X1 U15909 ( .B1(n14492), .B2(n14491), .A(n14490), .ZN(n14496) );
  XNOR2_X1 U15910 ( .A(n14493), .B(keyinput_56), .ZN(n14495) );
  XNOR2_X1 U15911 ( .A(P3_REG3_REG_20__SCAN_IN), .B(keyinput_55), .ZN(n14494)
         );
  NOR3_X1 U15912 ( .A1(n14496), .A2(n14495), .A3(n14494), .ZN(n14504) );
  XOR2_X1 U15913 ( .A(P3_REG3_REG_11__SCAN_IN), .B(keyinput_58), .Z(n14501) );
  XNOR2_X1 U15914 ( .A(n14497), .B(keyinput_57), .ZN(n14500) );
  XNOR2_X1 U15915 ( .A(P3_REG3_REG_18__SCAN_IN), .B(keyinput_60), .ZN(n14499)
         );
  XNOR2_X1 U15916 ( .A(P3_REG3_REG_2__SCAN_IN), .B(keyinput_59), .ZN(n14498)
         );
  NAND4_X1 U15917 ( .A1(n14501), .A2(n14500), .A3(n14499), .A4(n14498), .ZN(
        n14503) );
  XOR2_X1 U15918 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput_61), .Z(n14502) );
  OAI21_X1 U15919 ( .B1(n14504), .B2(n14503), .A(n14502), .ZN(n14508) );
  XNOR2_X1 U15920 ( .A(n14505), .B(keyinput_62), .ZN(n14507) );
  XNOR2_X1 U15921 ( .A(P3_REG3_REG_15__SCAN_IN), .B(keyinput_63), .ZN(n14506)
         );
  AOI21_X1 U15922 ( .B1(n14508), .B2(n14507), .A(n14506), .ZN(n14514) );
  XNOR2_X1 U15923 ( .A(P3_B_REG_SCAN_IN), .B(keyinput_64), .ZN(n14513) );
  XOR2_X1 U15924 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .Z(n14511)
         );
  XOR2_X1 U15925 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(keyinput_66), .Z(n14510)
         );
  XNOR2_X1 U15926 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .ZN(n14509)
         );
  NOR3_X1 U15927 ( .A1(n14511), .A2(n14510), .A3(n14509), .ZN(n14512) );
  OAI21_X1 U15928 ( .B1(n14514), .B2(n14513), .A(n14512), .ZN(n14517) );
  XOR2_X1 U15929 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .Z(n14516)
         );
  XNOR2_X1 U15930 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(keyinput_69), .ZN(n14515)
         );
  NAND3_X1 U15931 ( .A1(n14517), .A2(n14516), .A3(n14515), .ZN(n14520) );
  XOR2_X1 U15932 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(keyinput_70), .Z(n14519)
         );
  XOR2_X1 U15933 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .Z(n14518)
         );
  AOI21_X1 U15934 ( .B1(n14520), .B2(n14519), .A(n14518), .ZN(n14523) );
  XNOR2_X1 U15935 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .ZN(n14522)
         );
  XNOR2_X1 U15936 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .ZN(n14521)
         );
  NOR3_X1 U15937 ( .A1(n14523), .A2(n14522), .A3(n14521), .ZN(n14527) );
  XOR2_X1 U15938 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .Z(n14526)
         );
  XOR2_X1 U15939 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .Z(n14525)
         );
  XOR2_X1 U15940 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(keyinput_76), .Z(n14524)
         );
  OAI211_X1 U15941 ( .C1(n14527), .C2(n14526), .A(n14525), .B(n14524), .ZN(
        n14530) );
  XOR2_X1 U15942 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .Z(n14529)
         );
  XNOR2_X1 U15943 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .ZN(n14528)
         );
  NAND3_X1 U15944 ( .A1(n14530), .A2(n14529), .A3(n14528), .ZN(n14545) );
  INV_X1 U15945 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n14531) );
  OAI22_X1 U15946 ( .A1(keyinput_82), .A2(n14534), .B1(n14531), .B2(
        keyinput_83), .ZN(n14542) );
  OAI22_X1 U15947 ( .A1(n14533), .A2(keyinput_81), .B1(
        P3_DATAO_REG_11__SCAN_IN), .B2(keyinput_85), .ZN(n14541) );
  INV_X1 U15948 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n14532) );
  NOR2_X1 U15949 ( .A1(n14532), .A2(keyinput_79), .ZN(n14540) );
  AOI22_X1 U15950 ( .A1(n14532), .A2(keyinput_79), .B1(n14531), .B2(
        keyinput_83), .ZN(n14537) );
  AOI22_X1 U15951 ( .A1(P3_DATAO_REG_11__SCAN_IN), .A2(keyinput_85), .B1(
        P3_DATAO_REG_12__SCAN_IN), .B2(keyinput_84), .ZN(n14536) );
  AOI22_X1 U15952 ( .A1(n14534), .A2(keyinput_82), .B1(keyinput_81), .B2(
        n14533), .ZN(n14535) );
  AND3_X1 U15953 ( .A1(n14537), .A2(n14536), .A3(n14535), .ZN(n14538) );
  OAI21_X1 U15954 ( .B1(P3_DATAO_REG_12__SCAN_IN), .B2(keyinput_84), .A(n14538), .ZN(n14539) );
  NOR4_X1 U15955 ( .A1(n14542), .A2(n14541), .A3(n14540), .A4(n14539), .ZN(
        n14544) );
  XNOR2_X1 U15956 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(keyinput_80), .ZN(n14543)
         );
  NAND3_X1 U15957 ( .A1(n14545), .A2(n14544), .A3(n14543), .ZN(n14552) );
  XOR2_X1 U15958 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(keyinput_86), .Z(n14551)
         );
  XOR2_X1 U15959 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .Z(n14549) );
  XOR2_X1 U15960 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .Z(n14548) );
  XNOR2_X1 U15961 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(keyinput_87), .ZN(n14547)
         );
  XNOR2_X1 U15962 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(keyinput_90), .ZN(n14546)
         );
  NAND4_X1 U15963 ( .A1(n14549), .A2(n14548), .A3(n14547), .A4(n14546), .ZN(
        n14550) );
  AOI21_X1 U15964 ( .B1(n14552), .B2(n14551), .A(n14550), .ZN(n14559) );
  XOR2_X1 U15965 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(keyinput_91), .Z(n14555) );
  XNOR2_X1 U15966 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(keyinput_93), .ZN(n14554)
         );
  XNOR2_X1 U15967 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(keyinput_92), .ZN(n14553)
         );
  NAND3_X1 U15968 ( .A1(n14555), .A2(n14554), .A3(n14553), .ZN(n14558) );
  XOR2_X1 U15969 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(keyinput_94), .Z(n14557) );
  XNOR2_X1 U15970 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(keyinput_95), .ZN(n14556)
         );
  OAI211_X1 U15971 ( .C1(n14559), .C2(n14558), .A(n14557), .B(n14556), .ZN(
        n14565) );
  XOR2_X1 U15972 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(keyinput_96), .Z(n14564) );
  XNOR2_X1 U15973 ( .A(P3_ADDR_REG_0__SCAN_IN), .B(keyinput_97), .ZN(n14563)
         );
  INV_X1 U15974 ( .A(keyinput_100), .ZN(n14560) );
  XNOR2_X1 U15975 ( .A(n14560), .B(P3_ADDR_REG_3__SCAN_IN), .ZN(n14562) );
  XNOR2_X1 U15976 ( .A(P3_ADDR_REG_2__SCAN_IN), .B(keyinput_99), .ZN(n14561)
         );
  NAND2_X1 U15977 ( .A1(n14562), .A2(n14561), .ZN(n14568) );
  AOI211_X1 U15978 ( .C1(n14565), .C2(n14564), .A(n14563), .B(n14568), .ZN(
        n14572) );
  XOR2_X1 U15979 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(keyinput_98), .Z(n14567) );
  XOR2_X1 U15980 ( .A(P3_ADDR_REG_4__SCAN_IN), .B(keyinput_101), .Z(n14566) );
  OAI21_X1 U15981 ( .B1(n14568), .B2(n14567), .A(n14566), .ZN(n14571) );
  XOR2_X1 U15982 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(keyinput_103), .Z(n14570) );
  XNOR2_X1 U15983 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(keyinput_102), .ZN(n14569)
         );
  OAI211_X1 U15984 ( .C1(n14572), .C2(n14571), .A(n14570), .B(n14569), .ZN(
        n14575) );
  XOR2_X1 U15985 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(keyinput_104), .Z(n14574) );
  XOR2_X1 U15986 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(keyinput_105), .Z(n14573) );
  AOI21_X1 U15987 ( .B1(n14575), .B2(n14574), .A(n14573), .ZN(n14578) );
  XNOR2_X1 U15988 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(keyinput_106), .ZN(n14577)
         );
  XNOR2_X1 U15989 ( .A(n16160), .B(keyinput_107), .ZN(n14576) );
  OAI21_X1 U15990 ( .B1(n14578), .B2(n14577), .A(n14576), .ZN(n14582) );
  XNOR2_X1 U15991 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_108), .ZN(n14581) );
  XNOR2_X1 U15992 ( .A(n14579), .B(keyinput_109), .ZN(n14580) );
  AOI21_X1 U15993 ( .B1(n14582), .B2(n14581), .A(n14580), .ZN(n14586) );
  XOR2_X1 U15994 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_110), .Z(n14585) );
  XNOR2_X1 U15995 ( .A(n14583), .B(keyinput_111), .ZN(n14584) );
  OAI21_X1 U15996 ( .B1(n14586), .B2(n14585), .A(n14584), .ZN(n14591) );
  XNOR2_X1 U15997 ( .A(n14587), .B(keyinput_113), .ZN(n14590) );
  XNOR2_X1 U15998 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_112), .ZN(n14589) );
  XNOR2_X1 U15999 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_114), .ZN(n14588) );
  NAND4_X1 U16000 ( .A1(n14591), .A2(n14590), .A3(n14589), .A4(n14588), .ZN(
        n14595) );
  XOR2_X1 U16001 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_115), .Z(n14594) );
  XNOR2_X1 U16002 ( .A(n14592), .B(keyinput_116), .ZN(n14593) );
  AOI21_X1 U16003 ( .B1(n14595), .B2(n14594), .A(n14593), .ZN(n14598) );
  XOR2_X1 U16004 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_117), .Z(n14597) );
  XNOR2_X1 U16005 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_118), .ZN(n14596)
         );
  OAI21_X1 U16006 ( .B1(n14598), .B2(n14597), .A(n14596), .ZN(n14605) );
  XOR2_X1 U16007 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_121), .Z(n14602) );
  XNOR2_X1 U16008 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_122), .ZN(n14601)
         );
  XNOR2_X1 U16009 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_119), .ZN(n14600)
         );
  XNOR2_X1 U16010 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_120), .ZN(n14599)
         );
  NOR4_X1 U16011 ( .A1(n14602), .A2(n14601), .A3(n14600), .A4(n14599), .ZN(
        n14604) );
  XNOR2_X1 U16012 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_123), .ZN(n14603)
         );
  AOI21_X1 U16013 ( .B1(n14605), .B2(n14604), .A(n14603), .ZN(n14612) );
  XNOR2_X1 U16014 ( .A(n14606), .B(keyinput_124), .ZN(n14610) );
  XNOR2_X1 U16015 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_125), .ZN(n14609)
         );
  XNOR2_X1 U16016 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_127), .ZN(n14608)
         );
  XNOR2_X1 U16017 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_126), .ZN(n14607)
         );
  NAND4_X1 U16018 ( .A1(n14610), .A2(n14609), .A3(n14608), .A4(n14607), .ZN(
        n14611) );
  NOR3_X1 U16019 ( .A1(n14613), .A2(n14612), .A3(n14611), .ZN(n14614) );
  XOR2_X1 U16020 ( .A(n14615), .B(n14614), .Z(P2_U3194) );
  AOI21_X1 U16021 ( .B1(n14617), .B2(n14616), .A(n14686), .ZN(n14619) );
  NAND2_X1 U16022 ( .A1(n14619), .A2(n14618), .ZN(n14623) );
  AOI22_X1 U16023 ( .A1(n14700), .A2(n14934), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14622) );
  AOI22_X1 U16024 ( .A1(n14701), .A2(n14716), .B1(n14702), .B2(n14715), .ZN(
        n14621) );
  NAND2_X1 U16025 ( .A1(n15048), .A2(n14691), .ZN(n14620) );
  NAND4_X1 U16026 ( .A1(n14623), .A2(n14622), .A3(n14621), .A4(n14620), .ZN(
        P2_U3195) );
  INV_X1 U16027 ( .A(n14624), .ZN(n14625) );
  OAI21_X1 U16028 ( .B1(n14627), .B2(n14626), .A(n14625), .ZN(n14628) );
  XNOR2_X1 U16029 ( .A(n14629), .B(n14628), .ZN(n14630) );
  NAND2_X1 U16030 ( .A1(n14630), .A2(n14707), .ZN(n14637) );
  INV_X1 U16031 ( .A(n14631), .ZN(n14633) );
  NAND2_X1 U16032 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n16137)
         );
  INV_X1 U16033 ( .A(n16137), .ZN(n14632) );
  AOI21_X1 U16034 ( .B1(n14700), .B2(n14633), .A(n14632), .ZN(n14636) );
  AOI22_X1 U16035 ( .A1(n14701), .A2(n14725), .B1(n14702), .B2(n14723), .ZN(
        n14635) );
  NAND2_X1 U16036 ( .A1(n16606), .A2(n14691), .ZN(n14634) );
  NAND4_X1 U16037 ( .A1(n14637), .A2(n14636), .A3(n14635), .A4(n14634), .ZN(
        P2_U3196) );
  INV_X1 U16038 ( .A(n14638), .ZN(n14639) );
  AOI21_X1 U16039 ( .B1(n14652), .B2(n14639), .A(n14686), .ZN(n14642) );
  NOR3_X1 U16040 ( .A1(n14640), .A2(n14870), .A3(n14694), .ZN(n14641) );
  OAI21_X1 U16041 ( .B1(n14642), .B2(n14641), .A(n14693), .ZN(n14647) );
  INV_X1 U16042 ( .A(n14643), .ZN(n14875) );
  AOI22_X1 U16043 ( .A1(n14875), .A2(n14700), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14646) );
  AOI22_X1 U16044 ( .A1(n14838), .A2(n14702), .B1(n14701), .B2(n14714), .ZN(
        n14645) );
  NAND2_X1 U16045 ( .A1(n7953), .A2(n14691), .ZN(n14644) );
  NAND4_X1 U16046 ( .A1(n14647), .A2(n14646), .A3(n14645), .A4(n14644), .ZN(
        P2_U3197) );
  OAI22_X1 U16047 ( .A1(n14695), .A2(n14953), .B1(n14648), .B2(n14951), .ZN(
        n14882) );
  INV_X1 U16048 ( .A(n14882), .ZN(n14651) );
  AOI22_X1 U16049 ( .A1(n14700), .A2(n14887), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14649) );
  OAI21_X1 U16050 ( .B1(n14651), .B2(n14650), .A(n14649), .ZN(n14657) );
  INV_X1 U16051 ( .A(n14652), .ZN(n14653) );
  AOI211_X1 U16052 ( .C1(n14655), .C2(n14654), .A(n14686), .B(n14653), .ZN(
        n14656) );
  AOI211_X1 U16053 ( .C1(n15030), .C2(n14691), .A(n14657), .B(n14656), .ZN(
        n14658) );
  INV_X1 U16054 ( .A(n14658), .ZN(P2_U3201) );
  OAI21_X1 U16055 ( .B1(n14660), .B2(n14662), .A(n14659), .ZN(n14669) );
  NOR3_X1 U16056 ( .A1(n14662), .A2(n14661), .A3(n14694), .ZN(n14663) );
  OAI21_X1 U16057 ( .B1(n14663), .B2(n14701), .A(n14717), .ZN(n14667) );
  OAI22_X1 U16058 ( .A1(n14683), .A2(n14957), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14664), .ZN(n14665) );
  AOI21_X1 U16059 ( .B1(n14702), .B2(n14912), .A(n14665), .ZN(n14666) );
  OAI211_X1 U16060 ( .C1(n14960), .C2(n14705), .A(n14667), .B(n14666), .ZN(
        n14668) );
  AOI21_X1 U16061 ( .B1(n14707), .B2(n14669), .A(n14668), .ZN(n14670) );
  INV_X1 U16062 ( .A(n14670), .ZN(P2_U3205) );
  AOI22_X1 U16063 ( .A1(n14672), .A2(n14707), .B1(n14671), .B2(n14715), .ZN(
        n14679) );
  INV_X1 U16064 ( .A(n14673), .ZN(n14678) );
  AOI22_X1 U16065 ( .A1(n14701), .A2(n14912), .B1(n14702), .B2(n14914), .ZN(
        n14675) );
  NAND2_X1 U16066 ( .A1(P2_U3088), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n14674)
         );
  OAI211_X1 U16067 ( .C1(n14683), .C2(n14921), .A(n14675), .B(n14674), .ZN(
        n14676) );
  AOI21_X1 U16068 ( .B1(n15039), .B2(n14691), .A(n14676), .ZN(n14677) );
  OAI21_X1 U16069 ( .B1(n14679), .B2(n14678), .A(n14677), .ZN(P2_U3207) );
  OAI22_X1 U16070 ( .A1(n14950), .A2(n14953), .B1(n14680), .B2(n14951), .ZN(
        n14980) );
  AOI22_X1 U16071 ( .A1(n14681), .A2(n14980), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14682) );
  OAI21_X1 U16072 ( .B1(n14990), .B2(n14683), .A(n14682), .ZN(n14690) );
  INV_X1 U16073 ( .A(n14684), .ZN(n14685) );
  AOI211_X1 U16074 ( .C1(n14688), .C2(n14687), .A(n14686), .B(n14685), .ZN(
        n14689) );
  AOI211_X1 U16075 ( .C1(n15062), .C2(n14691), .A(n14690), .B(n14689), .ZN(
        n14692) );
  INV_X1 U16076 ( .A(n14692), .ZN(P2_U3210) );
  INV_X1 U16077 ( .A(n14693), .ZN(n14698) );
  NOR3_X1 U16078 ( .A1(n14696), .A2(n14695), .A3(n14694), .ZN(n14697) );
  AOI21_X1 U16079 ( .B1(n14698), .B2(n14707), .A(n14697), .ZN(n14711) );
  INV_X1 U16080 ( .A(n14699), .ZN(n14708) );
  AOI22_X1 U16081 ( .A1(n14854), .A2(n14700), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14704) );
  AOI22_X1 U16082 ( .A1(n14861), .A2(n14702), .B1(n14701), .B2(n14860), .ZN(
        n14703) );
  OAI211_X1 U16083 ( .C1(n14856), .C2(n14705), .A(n14704), .B(n14703), .ZN(
        n14706) );
  AOI21_X1 U16084 ( .B1(n14708), .B2(n14707), .A(n14706), .ZN(n14709) );
  OAI21_X1 U16085 ( .B1(n14711), .B2(n14710), .A(n14709), .ZN(P2_U3212) );
  MUX2_X1 U16086 ( .A(n14807), .B(P2_DATAO_REG_31__SCAN_IN), .S(n14736), .Z(
        P2_U3562) );
  MUX2_X1 U16087 ( .A(n14712), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14736), .Z(
        P2_U3561) );
  MUX2_X1 U16088 ( .A(n14713), .B(P2_DATAO_REG_29__SCAN_IN), .S(n14736), .Z(
        P2_U3560) );
  MUX2_X1 U16089 ( .A(n14839), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14736), .Z(
        P2_U3559) );
  MUX2_X1 U16090 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n14861), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U16091 ( .A(n14838), .B(P2_DATAO_REG_26__SCAN_IN), .S(n14736), .Z(
        P2_U3557) );
  MUX2_X1 U16092 ( .A(n14860), .B(P2_DATAO_REG_25__SCAN_IN), .S(n14736), .Z(
        P2_U3556) );
  MUX2_X1 U16093 ( .A(n14714), .B(P2_DATAO_REG_24__SCAN_IN), .S(n14736), .Z(
        P2_U3555) );
  MUX2_X1 U16094 ( .A(n14914), .B(P2_DATAO_REG_23__SCAN_IN), .S(n14736), .Z(
        P2_U3554) );
  MUX2_X1 U16095 ( .A(n14715), .B(P2_DATAO_REG_22__SCAN_IN), .S(n14736), .Z(
        P2_U3553) );
  MUX2_X1 U16096 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n14912), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U16097 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n14716), .S(P2_U3947), .Z(
        P2_U3551) );
  MUX2_X1 U16098 ( .A(n14717), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14736), .Z(
        P2_U3550) );
  MUX2_X1 U16099 ( .A(n14718), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14736), .Z(
        P2_U3549) );
  MUX2_X1 U16100 ( .A(n14719), .B(P2_DATAO_REG_17__SCAN_IN), .S(n14736), .Z(
        P2_U3548) );
  MUX2_X1 U16101 ( .A(n14720), .B(P2_DATAO_REG_16__SCAN_IN), .S(n14736), .Z(
        P2_U3547) );
  MUX2_X1 U16102 ( .A(n14721), .B(P2_DATAO_REG_15__SCAN_IN), .S(n14736), .Z(
        P2_U3546) );
  MUX2_X1 U16103 ( .A(n14722), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14736), .Z(
        P2_U3545) );
  MUX2_X1 U16104 ( .A(n14723), .B(P2_DATAO_REG_13__SCAN_IN), .S(n14736), .Z(
        P2_U3544) );
  MUX2_X1 U16105 ( .A(n14724), .B(P2_DATAO_REG_12__SCAN_IN), .S(n14736), .Z(
        P2_U3543) );
  MUX2_X1 U16106 ( .A(n14725), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14736), .Z(
        P2_U3542) );
  MUX2_X1 U16107 ( .A(n14726), .B(P2_DATAO_REG_10__SCAN_IN), .S(n14736), .Z(
        P2_U3541) );
  MUX2_X1 U16108 ( .A(n14727), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14736), .Z(
        P2_U3540) );
  MUX2_X1 U16109 ( .A(n14728), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14736), .Z(
        P2_U3539) );
  MUX2_X1 U16110 ( .A(n14729), .B(P2_DATAO_REG_7__SCAN_IN), .S(n14736), .Z(
        P2_U3538) );
  MUX2_X1 U16111 ( .A(n14730), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14736), .Z(
        P2_U3537) );
  MUX2_X1 U16112 ( .A(n14731), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14736), .Z(
        P2_U3536) );
  MUX2_X1 U16113 ( .A(n14732), .B(P2_DATAO_REG_4__SCAN_IN), .S(n14736), .Z(
        P2_U3535) );
  MUX2_X1 U16114 ( .A(n14733), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14736), .Z(
        P2_U3534) );
  MUX2_X1 U16115 ( .A(n14734), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14736), .Z(
        P2_U3533) );
  MUX2_X1 U16116 ( .A(n14735), .B(P2_DATAO_REG_1__SCAN_IN), .S(n14736), .Z(
        P2_U3532) );
  MUX2_X1 U16117 ( .A(n14737), .B(P2_DATAO_REG_0__SCAN_IN), .S(n14736), .Z(
        P2_U3531) );
  OAI211_X1 U16118 ( .C1(n14740), .C2(n14739), .A(n16152), .B(n14738), .ZN(
        n14749) );
  OAI211_X1 U16119 ( .C1(n14743), .C2(n14742), .A(n16148), .B(n14741), .ZN(
        n14748) );
  AND2_X1 U16120 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n14744) );
  AOI21_X1 U16121 ( .B1(n16110), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n14744), .ZN(
        n14747) );
  INV_X1 U16122 ( .A(n16127), .ZN(n16150) );
  NAND2_X1 U16123 ( .A1(n16150), .A2(n14745), .ZN(n14746) );
  NAND4_X1 U16124 ( .A1(n14749), .A2(n14748), .A3(n14747), .A4(n14746), .ZN(
        P2_U3217) );
  OAI211_X1 U16125 ( .C1(n14752), .C2(n14751), .A(n16152), .B(n14750), .ZN(
        n14761) );
  MUX2_X1 U16126 ( .A(n10289), .B(P2_REG1_REG_5__SCAN_IN), .S(n14756), .Z(
        n14753) );
  NAND3_X1 U16127 ( .A1(n16072), .A2(n14754), .A3(n14753), .ZN(n14755) );
  NAND3_X1 U16128 ( .A1(n16148), .A2(n14767), .A3(n14755), .ZN(n14760) );
  NAND2_X1 U16129 ( .A1(n16150), .A2(n14756), .ZN(n14759) );
  AND2_X1 U16130 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n14757) );
  AOI21_X1 U16131 ( .B1(n16110), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n14757), .ZN(
        n14758) );
  NAND4_X1 U16132 ( .A1(n14761), .A2(n14760), .A3(n14759), .A4(n14758), .ZN(
        P2_U3219) );
  OAI211_X1 U16133 ( .C1(n14764), .C2(n14763), .A(n16152), .B(n14762), .ZN(
        n14775) );
  MUX2_X1 U16134 ( .A(n10292), .B(P2_REG1_REG_6__SCAN_IN), .S(n14769), .Z(
        n14765) );
  NAND3_X1 U16135 ( .A1(n14767), .A2(n14766), .A3(n14765), .ZN(n14768) );
  NAND3_X1 U16136 ( .A1(n16148), .A2(n14781), .A3(n14768), .ZN(n14774) );
  NAND2_X1 U16137 ( .A1(n16150), .A2(n14769), .ZN(n14773) );
  INV_X1 U16138 ( .A(n14770), .ZN(n14771) );
  AOI21_X1 U16139 ( .B1(n16110), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n14771), .ZN(
        n14772) );
  NAND4_X1 U16140 ( .A1(n14775), .A2(n14774), .A3(n14773), .A4(n14772), .ZN(
        P2_U3220) );
  OAI211_X1 U16141 ( .C1(n14778), .C2(n14777), .A(n16152), .B(n14776), .ZN(
        n14789) );
  MUX2_X1 U16142 ( .A(n10295), .B(P2_REG1_REG_7__SCAN_IN), .S(n14783), .Z(
        n14779) );
  NAND3_X1 U16143 ( .A1(n14781), .A2(n14780), .A3(n14779), .ZN(n14782) );
  NAND3_X1 U16144 ( .A1(n16148), .A2(n14794), .A3(n14782), .ZN(n14788) );
  NAND2_X1 U16145 ( .A1(n16150), .A2(n14783), .ZN(n14787) );
  INV_X1 U16146 ( .A(n14784), .ZN(n14785) );
  AOI21_X1 U16147 ( .B1(n16110), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n14785), .ZN(
        n14786) );
  NAND4_X1 U16148 ( .A1(n14789), .A2(n14788), .A3(n14787), .A4(n14786), .ZN(
        P2_U3221) );
  OAI211_X1 U16149 ( .C1(n14791), .C2(n14790), .A(n16152), .B(n16140), .ZN(
        n14803) );
  MUX2_X1 U16150 ( .A(n10298), .B(P2_REG1_REG_8__SCAN_IN), .S(n14797), .Z(
        n14792) );
  NAND3_X1 U16151 ( .A1(n14794), .A2(n14793), .A3(n14792), .ZN(n14795) );
  NAND3_X1 U16152 ( .A1(n16148), .A2(n14796), .A3(n14795), .ZN(n14802) );
  NAND2_X1 U16153 ( .A1(n16150), .A2(n14797), .ZN(n14801) );
  INV_X1 U16154 ( .A(n14798), .ZN(n14799) );
  AOI21_X1 U16155 ( .B1(n16110), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n14799), .ZN(
        n14800) );
  NAND4_X1 U16156 ( .A1(n14803), .A2(n14802), .A3(n14801), .A4(n14800), .ZN(
        P2_U3222) );
  XNOR2_X1 U16157 ( .A(n14812), .B(n14804), .ZN(n14805) );
  NAND2_X1 U16158 ( .A1(n14805), .A2(n14930), .ZN(n14999) );
  NAND2_X1 U16159 ( .A1(n14807), .A2(n14806), .ZN(n15001) );
  NOR2_X1 U16160 ( .A1(n14992), .A2(n15001), .ZN(n14816) );
  NOR2_X1 U16161 ( .A1(n15000), .A2(n16515), .ZN(n14808) );
  AOI211_X1 U16162 ( .C1(n14992), .C2(P2_REG2_REG_31__SCAN_IN), .A(n14816), 
        .B(n14808), .ZN(n14809) );
  OAI21_X1 U16163 ( .B1(n14999), .B2(n14926), .A(n14809), .ZN(P2_U3234) );
  INV_X1 U16164 ( .A(n14811), .ZN(n14814) );
  OAI211_X1 U16165 ( .C1(n15003), .C2(n14814), .A(n14813), .B(n14930), .ZN(
        n15002) );
  NOR2_X1 U16166 ( .A1(n15003), .A2(n16515), .ZN(n14815) );
  AOI211_X1 U16167 ( .C1(n14992), .C2(P2_REG2_REG_30__SCAN_IN), .A(n14816), 
        .B(n14815), .ZN(n14817) );
  OAI21_X1 U16168 ( .B1(n14926), .B2(n15002), .A(n14817), .ZN(P2_U3235) );
  XNOR2_X1 U16169 ( .A(n14818), .B(n14822), .ZN(n14828) );
  OAI22_X1 U16170 ( .A1(n14820), .A2(n14953), .B1(n14819), .B2(n14951), .ZN(
        n14823) );
  AOI211_X1 U16171 ( .C1(n15011), .C2(n14844), .A(n14986), .B(n14824), .ZN(
        n15010) );
  AOI22_X1 U16172 ( .A1(n14825), .A2(n16511), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n14992), .ZN(n14826) );
  OAI21_X1 U16173 ( .B1(n14827), .B2(n16515), .A(n14826), .ZN(n14831) );
  INV_X1 U16174 ( .A(n14828), .ZN(n15014) );
  NOR2_X1 U16175 ( .A1(n15014), .A2(n14829), .ZN(n14830) );
  OAI21_X1 U16176 ( .B1(n15013), .B2(n14992), .A(n14832), .ZN(P2_U3237) );
  XNOR2_X1 U16177 ( .A(n14833), .B(n14834), .ZN(n15018) );
  NOR2_X1 U16178 ( .A1(n14835), .A2(n14834), .ZN(n14836) );
  OAI21_X1 U16179 ( .B1(n14837), .B2(n14836), .A(n14981), .ZN(n14841) );
  AOI22_X1 U16180 ( .A1(n14839), .A2(n14913), .B1(n14911), .B2(n14838), .ZN(
        n14840) );
  NAND2_X1 U16181 ( .A1(n14841), .A2(n14840), .ZN(n14842) );
  AOI21_X1 U16182 ( .B1(n15018), .B2(n16507), .A(n14842), .ZN(n15020) );
  AOI21_X1 U16183 ( .B1(n14843), .B2(n14852), .A(n14986), .ZN(n14845) );
  NAND2_X1 U16184 ( .A1(n14845), .A2(n14844), .ZN(n15015) );
  NOR2_X1 U16185 ( .A1(n15015), .A2(n14926), .ZN(n14849) );
  AOI22_X1 U16186 ( .A1(n14846), .A2(n16511), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14992), .ZN(n14847) );
  OAI21_X1 U16187 ( .B1(n15016), .B2(n16515), .A(n14847), .ZN(n14848) );
  AOI211_X1 U16188 ( .C1(n15018), .C2(n16519), .A(n14849), .B(n14848), .ZN(
        n14850) );
  OAI21_X1 U16189 ( .B1(n15020), .B2(n14992), .A(n14850), .ZN(P2_U3238) );
  XNOR2_X1 U16190 ( .A(n14851), .B(n14859), .ZN(n15025) );
  INV_X1 U16191 ( .A(n14872), .ZN(n14853) );
  AOI211_X1 U16192 ( .C1(n15022), .C2(n14853), .A(n14873), .B(n7427), .ZN(
        n15021) );
  AOI22_X1 U16193 ( .A1(n14854), .A2(n16511), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14992), .ZN(n14855) );
  OAI21_X1 U16194 ( .B1(n14856), .B2(n16515), .A(n14855), .ZN(n14864) );
  OAI21_X1 U16195 ( .B1(n14859), .B2(n14858), .A(n14857), .ZN(n14862) );
  AOI222_X1 U16196 ( .A1(n14981), .A2(n14862), .B1(n14861), .B2(n14913), .C1(
        n14860), .C2(n14911), .ZN(n15024) );
  NOR2_X1 U16197 ( .A1(n15024), .A2(n14992), .ZN(n14863) );
  AOI211_X1 U16198 ( .C1(n15021), .C2(n16508), .A(n14864), .B(n14863), .ZN(
        n14865) );
  OAI21_X1 U16199 ( .B1(n14892), .B2(n15025), .A(n14865), .ZN(P2_U3239) );
  XNOR2_X1 U16200 ( .A(n14866), .B(n14868), .ZN(n15029) );
  XOR2_X1 U16201 ( .A(n14868), .B(n14867), .Z(n14869) );
  OAI222_X1 U16202 ( .A1(n14953), .A2(n14871), .B1(n14951), .B2(n14870), .C1(
        n14949), .C2(n14869), .ZN(n15026) );
  NAND2_X1 U16203 ( .A1(n15026), .A2(n14954), .ZN(n14880) );
  INV_X1 U16204 ( .A(n14885), .ZN(n14874) );
  AOI211_X1 U16205 ( .C1(n7953), .C2(n14874), .A(n14873), .B(n14872), .ZN(
        n15027) );
  AOI22_X1 U16206 ( .A1(n14875), .A2(n16511), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14992), .ZN(n14876) );
  OAI21_X1 U16207 ( .B1(n14877), .B2(n16515), .A(n14876), .ZN(n14878) );
  AOI21_X1 U16208 ( .B1(n15027), .B2(n16508), .A(n14878), .ZN(n14879) );
  OAI211_X1 U16209 ( .C1(n14892), .C2(n15029), .A(n14880), .B(n14879), .ZN(
        P2_U3240) );
  XNOR2_X1 U16210 ( .A(n14891), .B(n14881), .ZN(n14883) );
  AOI21_X1 U16211 ( .B1(n14883), .B2(n14981), .A(n14882), .ZN(n15032) );
  NOR2_X1 U16212 ( .A1(n14889), .A2(n14903), .ZN(n14886) );
  AOI22_X1 U16213 ( .A1(n14992), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n14887), 
        .B2(n16511), .ZN(n14888) );
  OAI21_X1 U16214 ( .B1(n14889), .B2(n16515), .A(n14888), .ZN(n14894) );
  AOI21_X1 U16215 ( .B1(n14891), .B2(n14890), .A(n7492), .ZN(n15033) );
  NOR2_X1 U16216 ( .A1(n15033), .A2(n14892), .ZN(n14893) );
  AOI211_X1 U16217 ( .C1(n8425), .C2(n16508), .A(n14894), .B(n14893), .ZN(
        n14895) );
  OAI21_X1 U16218 ( .B1(n14992), .B2(n15032), .A(n14895), .ZN(P2_U3241) );
  XNOR2_X1 U16219 ( .A(n14896), .B(n14900), .ZN(n14898) );
  AOI21_X1 U16220 ( .B1(n14898), .B2(n14981), .A(n14897), .ZN(n15037) );
  XOR2_X1 U16221 ( .A(n14900), .B(n14899), .Z(n15038) );
  INV_X1 U16222 ( .A(n15038), .ZN(n14908) );
  NAND2_X1 U16223 ( .A1(n15035), .A2(n14918), .ZN(n14901) );
  NAND2_X1 U16224 ( .A1(n14901), .A2(n14930), .ZN(n14902) );
  NOR2_X1 U16225 ( .A1(n14903), .A2(n14902), .ZN(n15034) );
  NAND2_X1 U16226 ( .A1(n15034), .A2(n16508), .ZN(n14906) );
  AOI22_X1 U16227 ( .A1(n14992), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n14904), 
        .B2(n16511), .ZN(n14905) );
  OAI211_X1 U16228 ( .C1(n7952), .C2(n16515), .A(n14906), .B(n14905), .ZN(
        n14907) );
  AOI21_X1 U16229 ( .B1(n14908), .B2(n16417), .A(n14907), .ZN(n14909) );
  OAI21_X1 U16230 ( .B1(n14992), .B2(n15037), .A(n14909), .ZN(P2_U3242) );
  OAI21_X1 U16231 ( .B1(n7770), .B2(n7520), .A(n14910), .ZN(n14915) );
  AOI222_X1 U16232 ( .A1(n14981), .A2(n14915), .B1(n14914), .B2(n14913), .C1(
        n14912), .C2(n14911), .ZN(n15045) );
  INV_X1 U16233 ( .A(n14933), .ZN(n14916) );
  AOI21_X1 U16234 ( .B1(n15039), .B2(n14916), .A(n14986), .ZN(n14917) );
  NAND2_X1 U16235 ( .A1(n14918), .A2(n14917), .ZN(n15042) );
  NAND2_X1 U16236 ( .A1(n14919), .A2(n7770), .ZN(n15040) );
  NAND3_X1 U16237 ( .A1(n15041), .A2(n15040), .A3(n16417), .ZN(n14925) );
  NAND2_X1 U16238 ( .A1(n14992), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n14920) );
  OAI21_X1 U16239 ( .B1(n14922), .B2(n14921), .A(n14920), .ZN(n14923) );
  AOI21_X1 U16240 ( .B1(n15039), .B2(n16419), .A(n14923), .ZN(n14924) );
  OAI211_X1 U16241 ( .C1(n15042), .C2(n14926), .A(n14925), .B(n14924), .ZN(
        n14927) );
  INV_X1 U16242 ( .A(n14927), .ZN(n14928) );
  OAI21_X1 U16243 ( .B1(n15045), .B2(n14992), .A(n14928), .ZN(P2_U3243) );
  XOR2_X1 U16244 ( .A(n14938), .B(n14929), .Z(n15050) );
  NAND2_X1 U16245 ( .A1(n14955), .A2(n15048), .ZN(n14931) );
  NAND2_X1 U16246 ( .A1(n14931), .A2(n14930), .ZN(n14932) );
  NOR2_X1 U16247 ( .A1(n14933), .A2(n14932), .ZN(n15047) );
  NAND2_X1 U16248 ( .A1(n15048), .A2(n16419), .ZN(n14936) );
  AOI22_X1 U16249 ( .A1(n14992), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n14934), 
        .B2(n16511), .ZN(n14935) );
  NAND2_X1 U16250 ( .A1(n14936), .A2(n14935), .ZN(n14937) );
  AOI21_X1 U16251 ( .B1(n15047), .B2(n16508), .A(n14937), .ZN(n14944) );
  XNOR2_X1 U16252 ( .A(n14939), .B(n14938), .ZN(n14940) );
  OAI222_X1 U16253 ( .A1(n14953), .A2(n14942), .B1(n14951), .B2(n14941), .C1(
        n14940), .C2(n14949), .ZN(n15046) );
  NAND2_X1 U16254 ( .A1(n15046), .A2(n14954), .ZN(n14943) );
  OAI211_X1 U16255 ( .C1(n15050), .C2(n14892), .A(n14944), .B(n14943), .ZN(
        P2_U3244) );
  XOR2_X1 U16256 ( .A(n14947), .B(n14945), .Z(n15055) );
  XOR2_X1 U16257 ( .A(n14947), .B(n14946), .Z(n14948) );
  OAI222_X1 U16258 ( .A1(n14953), .A2(n14952), .B1(n14951), .B2(n14950), .C1(
        n14949), .C2(n14948), .ZN(n15051) );
  NAND2_X1 U16259 ( .A1(n15051), .A2(n14954), .ZN(n14963) );
  INV_X1 U16260 ( .A(n14955), .ZN(n14956) );
  AOI211_X1 U16261 ( .C1(n15053), .C2(n14969), .A(n14986), .B(n14956), .ZN(
        n15052) );
  INV_X1 U16262 ( .A(n14957), .ZN(n14958) );
  AOI22_X1 U16263 ( .A1(n14992), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14958), 
        .B2(n16511), .ZN(n14959) );
  OAI21_X1 U16264 ( .B1(n14960), .B2(n16515), .A(n14959), .ZN(n14961) );
  AOI21_X1 U16265 ( .B1(n15052), .B2(n16508), .A(n14961), .ZN(n14962) );
  OAI211_X1 U16266 ( .C1(n15055), .C2(n14892), .A(n14963), .B(n14962), .ZN(
        P2_U3245) );
  XOR2_X1 U16267 ( .A(n14967), .B(n14964), .Z(n14966) );
  AOI21_X1 U16268 ( .B1(n14966), .B2(n14981), .A(n14965), .ZN(n15059) );
  OAI21_X1 U16269 ( .B1(n7426), .B2(n7583), .A(n14968), .ZN(n15060) );
  INV_X1 U16270 ( .A(n15060), .ZN(n14977) );
  AOI21_X1 U16271 ( .B1(n14989), .B2(n15057), .A(n14986), .ZN(n14970) );
  AND2_X1 U16272 ( .A1(n14970), .A2(n14969), .ZN(n15056) );
  NAND2_X1 U16273 ( .A1(n15056), .A2(n16508), .ZN(n14974) );
  INV_X1 U16274 ( .A(n14971), .ZN(n14972) );
  AOI22_X1 U16275 ( .A1(n14992), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14972), 
        .B2(n16511), .ZN(n14973) );
  OAI211_X1 U16276 ( .C1(n14975), .C2(n16515), .A(n14974), .B(n14973), .ZN(
        n14976) );
  AOI21_X1 U16277 ( .B1(n14977), .B2(n16417), .A(n14976), .ZN(n14978) );
  OAI21_X1 U16278 ( .B1(n14992), .B2(n15059), .A(n14978), .ZN(P2_U3246) );
  XNOR2_X1 U16279 ( .A(n14979), .B(n14984), .ZN(n14982) );
  AOI21_X1 U16280 ( .B1(n14982), .B2(n14981), .A(n14980), .ZN(n15064) );
  XOR2_X1 U16281 ( .A(n14983), .B(n14984), .Z(n15065) );
  INV_X1 U16282 ( .A(n15065), .ZN(n14997) );
  INV_X1 U16283 ( .A(n14985), .ZN(n14987) );
  AOI21_X1 U16284 ( .B1(n15062), .B2(n14987), .A(n14986), .ZN(n14988) );
  AND2_X1 U16285 ( .A1(n14989), .A2(n14988), .ZN(n15061) );
  NAND2_X1 U16286 ( .A1(n15061), .A2(n16508), .ZN(n14994) );
  INV_X1 U16287 ( .A(n14990), .ZN(n14991) );
  AOI22_X1 U16288 ( .A1(n14992), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14991), 
        .B2(n16511), .ZN(n14993) );
  OAI211_X1 U16289 ( .C1(n14995), .C2(n16515), .A(n14994), .B(n14993), .ZN(
        n14996) );
  AOI21_X1 U16290 ( .B1(n14997), .B2(n16417), .A(n14996), .ZN(n14998) );
  OAI21_X1 U16291 ( .B1(n16522), .B2(n15064), .A(n14998), .ZN(P2_U3247) );
  OAI211_X1 U16292 ( .C1(n15000), .C2(n16616), .A(n14999), .B(n15001), .ZN(
        n15086) );
  MUX2_X1 U16293 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n15086), .S(n7433), .Z(
        P2_U3530) );
  OAI211_X1 U16294 ( .C1(n15003), .C2(n16616), .A(n15002), .B(n15001), .ZN(
        n15087) );
  MUX2_X1 U16295 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n15087), .S(n7433), .Z(
        P2_U3529) );
  NAND2_X1 U16296 ( .A1(n15004), .A2(n16621), .ZN(n15008) );
  NAND2_X1 U16297 ( .A1(n15005), .A2(n15079), .ZN(n15007) );
  NAND4_X1 U16298 ( .A1(n15008), .A2(n15009), .A3(n15007), .A4(n15006), .ZN(
        n15088) );
  MUX2_X1 U16299 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n15088), .S(n7433), .Z(
        P2_U3528) );
  AOI21_X1 U16300 ( .B1(n15079), .B2(n15011), .A(n15010), .ZN(n15012) );
  OAI211_X1 U16301 ( .C1(n10450), .C2(n15014), .A(n15013), .B(n15012), .ZN(
        n15089) );
  MUX2_X1 U16302 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n15089), .S(n7433), .Z(
        P2_U3527) );
  OAI21_X1 U16303 ( .B1(n15016), .B2(n16616), .A(n15015), .ZN(n15017) );
  AOI21_X1 U16304 ( .B1(n15018), .B2(n16610), .A(n15017), .ZN(n15019) );
  NAND2_X1 U16305 ( .A1(n15020), .A2(n15019), .ZN(n15090) );
  MUX2_X1 U16306 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n15090), .S(n7433), .Z(
        P2_U3526) );
  AOI21_X1 U16307 ( .B1(n15079), .B2(n15022), .A(n15021), .ZN(n15023) );
  OAI211_X1 U16308 ( .C1(n15082), .C2(n15025), .A(n15024), .B(n15023), .ZN(
        n15091) );
  MUX2_X1 U16309 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n15091), .S(n7433), .Z(
        P2_U3525) );
  AOI211_X1 U16310 ( .C1(n15079), .C2(n7953), .A(n15027), .B(n15026), .ZN(
        n15028) );
  OAI21_X1 U16311 ( .B1(n15082), .B2(n15029), .A(n15028), .ZN(n15092) );
  MUX2_X1 U16312 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n15092), .S(n7433), .Z(
        P2_U3524) );
  AOI21_X1 U16313 ( .B1(n15079), .B2(n15030), .A(n8425), .ZN(n15031) );
  OAI211_X1 U16314 ( .C1(n15033), .C2(n15082), .A(n15032), .B(n15031), .ZN(
        n15093) );
  MUX2_X1 U16315 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n15093), .S(n7433), .Z(
        P2_U3523) );
  AOI21_X1 U16316 ( .B1(n15079), .B2(n15035), .A(n15034), .ZN(n15036) );
  OAI211_X1 U16317 ( .C1(n15038), .C2(n15082), .A(n15037), .B(n15036), .ZN(
        n15094) );
  MUX2_X1 U16318 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n15094), .S(n7433), .Z(
        P2_U3522) );
  NAND2_X1 U16319 ( .A1(n15039), .A2(n15079), .ZN(n15044) );
  NAND3_X1 U16320 ( .A1(n15041), .A2(n16621), .A3(n15040), .ZN(n15043) );
  NAND4_X1 U16321 ( .A1(n15045), .A2(n15044), .A3(n15043), .A4(n15042), .ZN(
        n15095) );
  MUX2_X1 U16322 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n15095), .S(n7433), .Z(
        P2_U3521) );
  AOI211_X1 U16323 ( .C1(n15079), .C2(n15048), .A(n15047), .B(n15046), .ZN(
        n15049) );
  OAI21_X1 U16324 ( .B1(n15082), .B2(n15050), .A(n15049), .ZN(n15096) );
  MUX2_X1 U16325 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n15096), .S(n7433), .Z(
        P2_U3520) );
  AOI211_X1 U16326 ( .C1(n15079), .C2(n15053), .A(n15052), .B(n15051), .ZN(
        n15054) );
  OAI21_X1 U16327 ( .B1(n15082), .B2(n15055), .A(n15054), .ZN(n15097) );
  MUX2_X1 U16328 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n15097), .S(n7433), .Z(
        P2_U3519) );
  AOI21_X1 U16329 ( .B1(n15079), .B2(n15057), .A(n15056), .ZN(n15058) );
  OAI211_X1 U16330 ( .C1(n15060), .C2(n15082), .A(n15059), .B(n15058), .ZN(
        n15098) );
  MUX2_X1 U16331 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n15098), .S(n7433), .Z(
        P2_U3518) );
  AOI21_X1 U16332 ( .B1(n15079), .B2(n15062), .A(n15061), .ZN(n15063) );
  OAI211_X1 U16333 ( .C1(n15065), .C2(n15082), .A(n15064), .B(n15063), .ZN(
        n15099) );
  MUX2_X1 U16334 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n15099), .S(n7433), .Z(
        P2_U3517) );
  INV_X1 U16335 ( .A(n15066), .ZN(n15071) );
  AOI21_X1 U16336 ( .B1(n15079), .B2(n15068), .A(n15067), .ZN(n15069) );
  OAI211_X1 U16337 ( .C1(n15071), .C2(n15082), .A(n15070), .B(n15069), .ZN(
        n15100) );
  MUX2_X1 U16338 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n15100), .S(n7433), .Z(
        P2_U3516) );
  AOI21_X1 U16339 ( .B1(n15079), .B2(n15073), .A(n15072), .ZN(n15074) );
  OAI211_X1 U16340 ( .C1(n15076), .C2(n15082), .A(n15075), .B(n15074), .ZN(
        n15101) );
  MUX2_X1 U16341 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n15101), .S(n7433), .Z(
        P2_U3515) );
  AOI21_X1 U16342 ( .B1(n15079), .B2(n15078), .A(n15077), .ZN(n15080) );
  OAI211_X1 U16343 ( .C1(n15083), .C2(n15082), .A(n15081), .B(n15080), .ZN(
        n15103) );
  MUX2_X1 U16344 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n15103), .S(n7433), .Z(
        P2_U3514) );
  MUX2_X1 U16345 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n15084), .S(n7433), .Z(
        P2_U3503) );
  MUX2_X1 U16346 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n15085), .S(n7433), .Z(
        P2_U3500) );
  MUX2_X1 U16347 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n15086), .S(n15102), .Z(
        P2_U3498) );
  MUX2_X1 U16348 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n15087), .S(n15102), .Z(
        P2_U3497) );
  MUX2_X1 U16349 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n15088), .S(n15102), .Z(
        P2_U3496) );
  MUX2_X1 U16350 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n15089), .S(n15102), .Z(
        P2_U3495) );
  MUX2_X1 U16351 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n15090), .S(n15102), .Z(
        P2_U3494) );
  MUX2_X1 U16352 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n15091), .S(n15102), .Z(
        P2_U3493) );
  MUX2_X1 U16353 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n15092), .S(n15102), .Z(
        P2_U3492) );
  MUX2_X1 U16354 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n15093), .S(n15102), .Z(
        P2_U3491) );
  MUX2_X1 U16355 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n15094), .S(n15102), .Z(
        P2_U3490) );
  MUX2_X1 U16356 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n15095), .S(n15102), .Z(
        P2_U3489) );
  MUX2_X1 U16357 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n15096), .S(n15102), .Z(
        P2_U3488) );
  MUX2_X1 U16358 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n15097), .S(n15102), .Z(
        P2_U3487) );
  MUX2_X1 U16359 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n15098), .S(n15102), .Z(
        P2_U3486) );
  MUX2_X1 U16360 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n15099), .S(n15102), .Z(
        P2_U3484) );
  MUX2_X1 U16361 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n15100), .S(n15102), .Z(
        P2_U3481) );
  MUX2_X1 U16362 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n15101), .S(n15102), .Z(
        P2_U3478) );
  MUX2_X1 U16363 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n15103), .S(n15102), .Z(
        P2_U3475) );
  INV_X1 U16364 ( .A(n15104), .ZN(n15973) );
  INV_X1 U16365 ( .A(n15105), .ZN(n15109) );
  NAND3_X1 U16366 ( .A1(n15106), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n15108) );
  OAI22_X1 U16367 ( .A1(n15109), .A2(n15108), .B1(n15107), .B2(n15133), .ZN(
        n15110) );
  INV_X1 U16368 ( .A(n15110), .ZN(n15111) );
  OAI21_X1 U16369 ( .B1(n15973), .B2(n15123), .A(n15111), .ZN(P2_U3296) );
  INV_X1 U16370 ( .A(n15112), .ZN(n15978) );
  OAI222_X1 U16371 ( .A1(n15131), .A2(n15978), .B1(n15114), .B2(P2_U3088), 
        .C1(n15113), .C2(n15133), .ZN(P2_U3298) );
  OAI222_X1 U16372 ( .A1(n15133), .A2(n15117), .B1(n15131), .B2(n15116), .C1(
        P2_U3088), .C2(n15115), .ZN(P2_U3299) );
  INV_X1 U16373 ( .A(n15118), .ZN(n15981) );
  OAI222_X1 U16374 ( .A1(n15133), .A2(n15120), .B1(n15123), .B2(n15981), .C1(
        P2_U3088), .C2(n15119), .ZN(P2_U3300) );
  INV_X1 U16375 ( .A(n15121), .ZN(n15124) );
  INV_X1 U16376 ( .A(n15122), .ZN(n15984) );
  OAI222_X1 U16377 ( .A1(n15133), .A2(n15125), .B1(n15124), .B2(P2_U3088), 
        .C1(n15123), .C2(n15984), .ZN(P2_U3301) );
  INV_X1 U16378 ( .A(n15126), .ZN(n15989) );
  OAI222_X1 U16379 ( .A1(n15133), .A2(n15128), .B1(n15131), .B2(n15989), .C1(
        P2_U3088), .C2(n15127), .ZN(P2_U3302) );
  INV_X1 U16380 ( .A(n15129), .ZN(n15994) );
  OAI222_X1 U16381 ( .A1(n15133), .A2(n15132), .B1(n15131), .B2(n15994), .C1(
        P2_U3088), .C2(n15130), .ZN(P2_U3303) );
  INV_X1 U16382 ( .A(n15134), .ZN(n15135) );
  MUX2_X1 U16383 ( .A(n15135), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI22_X1 U16384 ( .A1(n15621), .A2(n15136), .B1(n15636), .B2(n7462), .ZN(
        n15137) );
  XNOR2_X1 U16385 ( .A(n15137), .B(n15253), .ZN(n15139) );
  OAI22_X1 U16386 ( .A1(n15621), .A2(n7462), .B1(n15636), .B2(n15223), .ZN(
        n15138) );
  NOR2_X1 U16387 ( .A1(n15139), .A2(n15138), .ZN(n15250) );
  AOI21_X1 U16388 ( .B1(n15139), .B2(n15138), .A(n15250), .ZN(n15228) );
  AOI22_X1 U16389 ( .A1(n15883), .A2(n15255), .B1(n7432), .B2(n15736), .ZN(
        n15140) );
  XNOR2_X1 U16390 ( .A(n15140), .B(n15253), .ZN(n15187) );
  INV_X1 U16391 ( .A(n15187), .ZN(n15190) );
  AOI22_X1 U16392 ( .A1(n15883), .A2(n7432), .B1(n15252), .B2(n15736), .ZN(
        n15188) );
  INV_X1 U16393 ( .A(n15188), .ZN(n15189) );
  AND2_X1 U16394 ( .A1(n15550), .A2(n15252), .ZN(n15141) );
  AOI21_X1 U16395 ( .B1(n15889), .B2(n7432), .A(n15141), .ZN(n15184) );
  INV_X1 U16396 ( .A(n15184), .ZN(n15186) );
  NAND2_X1 U16397 ( .A1(n15889), .A2(n15255), .ZN(n15143) );
  NAND2_X1 U16398 ( .A1(n15550), .A2(n7432), .ZN(n15142) );
  NAND2_X1 U16399 ( .A1(n15143), .A2(n15142), .ZN(n15144) );
  XNOR2_X1 U16400 ( .A(n15144), .B(n15253), .ZN(n15185) );
  NAND2_X1 U16401 ( .A1(n15146), .A2(n15145), .ZN(n15147) );
  NAND2_X1 U16402 ( .A1(n15561), .A2(n15255), .ZN(n15150) );
  NAND2_X1 U16403 ( .A1(n15540), .A2(n7432), .ZN(n15149) );
  NAND2_X1 U16404 ( .A1(n15150), .A2(n15149), .ZN(n15151) );
  XNOR2_X1 U16405 ( .A(n15151), .B(n15253), .ZN(n15154) );
  AND2_X1 U16406 ( .A1(n15252), .A2(n15540), .ZN(n15152) );
  AOI21_X1 U16407 ( .B1(n15561), .B2(n7432), .A(n15152), .ZN(n15352) );
  NAND2_X1 U16408 ( .A1(n15353), .A2(n15352), .ZN(n15351) );
  INV_X1 U16409 ( .A(n15153), .ZN(n15156) );
  INV_X1 U16410 ( .A(n15154), .ZN(n15155) );
  NAND2_X1 U16411 ( .A1(n15156), .A2(n15155), .ZN(n15355) );
  NAND2_X1 U16412 ( .A1(n15919), .A2(n15255), .ZN(n15158) );
  NAND2_X1 U16413 ( .A1(n15788), .A2(n7432), .ZN(n15157) );
  NAND2_X1 U16414 ( .A1(n15158), .A2(n15157), .ZN(n15159) );
  XNOR2_X1 U16415 ( .A(n15159), .B(n15253), .ZN(n15160) );
  AOI22_X1 U16416 ( .A1(n15919), .A2(n7432), .B1(n15252), .B2(n15788), .ZN(
        n15161) );
  XNOR2_X1 U16417 ( .A(n15160), .B(n15161), .ZN(n15288) );
  INV_X1 U16418 ( .A(n15160), .ZN(n15162) );
  NAND2_X1 U16419 ( .A1(n15909), .A2(n15255), .ZN(n15164) );
  NAND2_X1 U16420 ( .A1(n15768), .A2(n7432), .ZN(n15163) );
  NAND2_X1 U16421 ( .A1(n15164), .A2(n15163), .ZN(n15165) );
  XNOR2_X1 U16422 ( .A(n15165), .B(n15221), .ZN(n15168) );
  AND2_X1 U16423 ( .A1(n15768), .A2(n15252), .ZN(n15166) );
  AOI21_X1 U16424 ( .B1(n15909), .B2(n7432), .A(n15166), .ZN(n15167) );
  NOR2_X1 U16425 ( .A1(n15168), .A2(n15167), .ZN(n15294) );
  NAND2_X1 U16426 ( .A1(n15778), .A2(n15255), .ZN(n15170) );
  NAND2_X1 U16427 ( .A1(n15790), .A2(n7432), .ZN(n15169) );
  NAND2_X1 U16428 ( .A1(n15170), .A2(n15169), .ZN(n15171) );
  XNOR2_X1 U16429 ( .A(n15171), .B(n15253), .ZN(n15175) );
  NAND2_X1 U16430 ( .A1(n15778), .A2(n7432), .ZN(n15173) );
  NAND2_X1 U16431 ( .A1(n15790), .A2(n15252), .ZN(n15172) );
  NAND2_X1 U16432 ( .A1(n15173), .A2(n15172), .ZN(n15174) );
  NOR2_X1 U16433 ( .A1(n15175), .A2(n15174), .ZN(n15176) );
  AOI21_X1 U16434 ( .B1(n15175), .B2(n15174), .A(n15176), .ZN(n15331) );
  NAND2_X1 U16435 ( .A1(n15746), .A2(n15255), .ZN(n15178) );
  NAND2_X1 U16436 ( .A1(n15769), .A2(n7432), .ZN(n15177) );
  NAND2_X1 U16437 ( .A1(n15178), .A2(n15177), .ZN(n15179) );
  XNOR2_X1 U16438 ( .A(n15179), .B(n15253), .ZN(n15182) );
  AOI22_X1 U16439 ( .A1(n15746), .A2(n7432), .B1(n15252), .B2(n15769), .ZN(
        n15180) );
  XNOR2_X1 U16440 ( .A(n15182), .B(n15180), .ZN(n15243) );
  INV_X1 U16441 ( .A(n15180), .ZN(n15181) );
  OR2_X1 U16442 ( .A1(n15182), .A2(n15181), .ZN(n15183) );
  XOR2_X1 U16443 ( .A(n15184), .B(n15185), .Z(n15311) );
  XOR2_X1 U16444 ( .A(n15188), .B(n15187), .Z(n15271) );
  OAI21_X1 U16445 ( .B1(n15190), .B2(n15189), .A(n15269), .ZN(n15319) );
  NAND2_X1 U16446 ( .A1(n15698), .A2(n15255), .ZN(n15192) );
  NAND2_X1 U16447 ( .A1(n15554), .A2(n7432), .ZN(n15191) );
  NAND2_X1 U16448 ( .A1(n15192), .A2(n15191), .ZN(n15193) );
  XNOR2_X1 U16449 ( .A(n15193), .B(n15253), .ZN(n15196) );
  NAND2_X1 U16450 ( .A1(n15698), .A2(n7432), .ZN(n15195) );
  NAND2_X1 U16451 ( .A1(n15554), .A2(n15252), .ZN(n15194) );
  NAND2_X1 U16452 ( .A1(n15195), .A2(n15194), .ZN(n15197) );
  NAND2_X1 U16453 ( .A1(n15196), .A2(n15197), .ZN(n15320) );
  INV_X1 U16454 ( .A(n15196), .ZN(n15199) );
  INV_X1 U16455 ( .A(n15197), .ZN(n15198) );
  NAND2_X1 U16456 ( .A1(n15199), .A2(n15198), .ZN(n15322) );
  NAND2_X1 U16457 ( .A1(n15318), .A2(n15322), .ZN(n15234) );
  INV_X1 U16458 ( .A(n15703), .ZN(n15557) );
  OAI22_X1 U16459 ( .A1(n15686), .A2(n7462), .B1(n15557), .B2(n15223), .ZN(
        n15204) );
  NAND2_X1 U16460 ( .A1(n15867), .A2(n15255), .ZN(n15201) );
  NAND2_X1 U16461 ( .A1(n15703), .A2(n7432), .ZN(n15200) );
  NAND2_X1 U16462 ( .A1(n15201), .A2(n15200), .ZN(n15202) );
  XNOR2_X1 U16463 ( .A(n15202), .B(n15253), .ZN(n15203) );
  XOR2_X1 U16464 ( .A(n15204), .B(n15203), .Z(n15235) );
  INV_X1 U16465 ( .A(n15203), .ZN(n15206) );
  INV_X1 U16466 ( .A(n15204), .ZN(n15205) );
  NAND2_X1 U16467 ( .A1(n15859), .A2(n15255), .ZN(n15208) );
  NAND2_X1 U16468 ( .A1(n15577), .A2(n7432), .ZN(n15207) );
  NAND2_X1 U16469 ( .A1(n15208), .A2(n15207), .ZN(n15209) );
  XNOR2_X1 U16470 ( .A(n15209), .B(n15253), .ZN(n15211) );
  INV_X1 U16471 ( .A(n15859), .ZN(n15578) );
  INV_X1 U16472 ( .A(n15577), .ZN(n15652) );
  OAI22_X1 U16473 ( .A1(n15578), .A2(n7462), .B1(n15652), .B2(n15223), .ZN(
        n15210) );
  XNOR2_X1 U16474 ( .A(n15211), .B(n15210), .ZN(n15303) );
  INV_X1 U16475 ( .A(n15853), .ZN(n15655) );
  INV_X1 U16476 ( .A(n15667), .ZN(n15579) );
  OAI22_X1 U16477 ( .A1(n15655), .A2(n7462), .B1(n15579), .B2(n15223), .ZN(
        n15216) );
  NAND2_X1 U16478 ( .A1(n15853), .A2(n15255), .ZN(n15213) );
  NAND2_X1 U16479 ( .A1(n15667), .A2(n7432), .ZN(n15212) );
  NAND2_X1 U16480 ( .A1(n15213), .A2(n15212), .ZN(n15214) );
  XNOR2_X1 U16481 ( .A(n15214), .B(n15253), .ZN(n15215) );
  XOR2_X1 U16482 ( .A(n15216), .B(n15215), .Z(n15281) );
  INV_X1 U16483 ( .A(n15215), .ZN(n15218) );
  INV_X1 U16484 ( .A(n15216), .ZN(n15217) );
  NAND2_X1 U16485 ( .A1(n15847), .A2(n15255), .ZN(n15220) );
  NAND2_X1 U16486 ( .A1(n15614), .A2(n7432), .ZN(n15219) );
  NAND2_X1 U16487 ( .A1(n15220), .A2(n15219), .ZN(n15222) );
  XNOR2_X1 U16488 ( .A(n15222), .B(n15221), .ZN(n15226) );
  NOR2_X1 U16489 ( .A1(n15653), .A2(n15223), .ZN(n15224) );
  AOI21_X1 U16490 ( .B1(n15847), .B2(n7432), .A(n15224), .ZN(n15225) );
  NOR2_X1 U16491 ( .A1(n15226), .A2(n15225), .ZN(n15343) );
  NAND2_X1 U16492 ( .A1(n15226), .A2(n15225), .ZN(n15341) );
  OAI21_X1 U16493 ( .B1(n15228), .B2(n15227), .A(n15251), .ZN(n15229) );
  NAND2_X1 U16494 ( .A1(n15229), .A2(n15332), .ZN(n15233) );
  NOR2_X1 U16495 ( .A1(n15359), .A2(n15653), .ZN(n15231) );
  INV_X1 U16496 ( .A(n15613), .ZN(n15581) );
  OAI22_X1 U16497 ( .A1(n15362), .A2(n15581), .B1(n15618), .B2(n15360), .ZN(
        n15230) );
  AOI211_X1 U16498 ( .C1(P1_REG3_REG_27__SCAN_IN), .C2(P1_U3086), .A(n15231), 
        .B(n15230), .ZN(n15232) );
  OAI211_X1 U16499 ( .C1(n15621), .C2(n15340), .A(n15233), .B(n15232), .ZN(
        P1_U3214) );
  XOR2_X1 U16500 ( .A(n15235), .B(n15234), .Z(n15240) );
  AND2_X1 U16501 ( .A1(n15789), .A2(n15577), .ZN(n15236) );
  AOI21_X1 U16502 ( .B1(n15554), .B2(n15787), .A(n15236), .ZN(n15682) );
  AOI22_X1 U16503 ( .A1(n15684), .A2(n15312), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15237) );
  OAI21_X1 U16504 ( .B1(n15682), .B2(n15264), .A(n15237), .ZN(n15238) );
  AOI21_X1 U16505 ( .B1(n15867), .B2(n15365), .A(n15238), .ZN(n15239) );
  OAI21_X1 U16506 ( .B1(n15240), .B2(n15367), .A(n15239), .ZN(P1_U3216) );
  INV_X1 U16507 ( .A(n15746), .ZN(n15897) );
  OAI21_X1 U16508 ( .B1(n15243), .B2(n15242), .A(n15241), .ZN(n15244) );
  NAND2_X1 U16509 ( .A1(n15244), .A2(n15332), .ZN(n15249) );
  NAND2_X1 U16510 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n15522)
         );
  INV_X1 U16511 ( .A(n15522), .ZN(n15247) );
  INV_X1 U16512 ( .A(n15550), .ZN(n15754) );
  INV_X1 U16513 ( .A(n15758), .ZN(n15245) );
  OAI22_X1 U16514 ( .A1(n15754), .A2(n15362), .B1(n15245), .B2(n15360), .ZN(
        n15246) );
  AOI211_X1 U16515 ( .C1(n15337), .C2(n15790), .A(n15247), .B(n15246), .ZN(
        n15248) );
  OAI211_X1 U16516 ( .C1(n15897), .C2(n15340), .A(n15249), .B(n15248), .ZN(
        P1_U3219) );
  AOI22_X1 U16517 ( .A1(n15837), .A2(n7432), .B1(n15252), .B2(n15613), .ZN(
        n15254) );
  XNOR2_X1 U16518 ( .A(n15254), .B(n15253), .ZN(n15257) );
  AOI22_X1 U16519 ( .A1(n15837), .A2(n15255), .B1(n7432), .B2(n15613), .ZN(
        n15256) );
  XNOR2_X1 U16520 ( .A(n15257), .B(n15256), .ZN(n15258) );
  XNOR2_X1 U16521 ( .A(n15259), .B(n15258), .ZN(n15268) );
  NOR2_X1 U16522 ( .A1(n15360), .A2(n15603), .ZN(n15266) );
  OR2_X1 U16523 ( .A1(n15636), .A2(n15805), .ZN(n15262) );
  OR2_X1 U16524 ( .A1(n15260), .A2(n16389), .ZN(n15261) );
  AND2_X1 U16525 ( .A1(n15262), .A2(n15261), .ZN(n15599) );
  OAI22_X1 U16526 ( .A1(n15264), .A2(n15599), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15263), .ZN(n15265) );
  AOI211_X1 U16527 ( .C1(n15837), .C2(n15365), .A(n15266), .B(n15265), .ZN(
        n15267) );
  OAI21_X1 U16528 ( .B1(n15268), .B2(n15367), .A(n15267), .ZN(P1_U3220) );
  INV_X1 U16529 ( .A(n15883), .ZN(n15723) );
  OAI21_X1 U16530 ( .B1(n15271), .B2(n15270), .A(n15269), .ZN(n15272) );
  NAND2_X1 U16531 ( .A1(n15272), .A2(n15332), .ZN(n15279) );
  NAND2_X1 U16532 ( .A1(n15554), .A2(n15789), .ZN(n15274) );
  NAND2_X1 U16533 ( .A1(n15550), .A2(n15787), .ZN(n15273) );
  NAND2_X1 U16534 ( .A1(n15274), .A2(n15273), .ZN(n15715) );
  OAI22_X1 U16535 ( .A1(n15720), .A2(n15360), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15275), .ZN(n15276) );
  AOI21_X1 U16536 ( .B1(n15715), .B2(n15277), .A(n15276), .ZN(n15278) );
  OAI211_X1 U16537 ( .C1(n15723), .C2(n15340), .A(n15279), .B(n15278), .ZN(
        P1_U3223) );
  XOR2_X1 U16538 ( .A(n15281), .B(n15280), .Z(n15286) );
  INV_X1 U16539 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n15282) );
  OAI22_X1 U16540 ( .A1(n15362), .A2(n15653), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15282), .ZN(n15284) );
  OAI22_X1 U16541 ( .A1(n15359), .A2(n15652), .B1(n15360), .B2(n15656), .ZN(
        n15283) );
  AOI211_X1 U16542 ( .C1(n15853), .C2(n15365), .A(n15284), .B(n15283), .ZN(
        n15285) );
  OAI21_X1 U16543 ( .B1(n15286), .B2(n15367), .A(n15285), .ZN(P1_U3225) );
  XOR2_X1 U16544 ( .A(n15288), .B(n15287), .Z(n15293) );
  INV_X1 U16545 ( .A(n15540), .ZN(n15806) );
  OAI21_X1 U16546 ( .B1(n15359), .B2(n15806), .A(n15289), .ZN(n15291) );
  OAI22_X1 U16547 ( .A1(n15362), .A2(n15807), .B1(n15804), .B2(n15360), .ZN(
        n15290) );
  AOI211_X1 U16548 ( .C1(n15919), .C2(n15365), .A(n15291), .B(n15290), .ZN(
        n15292) );
  OAI21_X1 U16549 ( .B1(n15293), .B2(n15367), .A(n15292), .ZN(P1_U3226) );
  NOR2_X1 U16550 ( .A1(n15294), .A2(n7562), .ZN(n15295) );
  XNOR2_X1 U16551 ( .A(n15296), .B(n15295), .ZN(n15301) );
  INV_X1 U16552 ( .A(n15788), .ZN(n15564) );
  OAI21_X1 U16553 ( .B1(n15359), .B2(n15564), .A(n15297), .ZN(n15299) );
  OAI22_X1 U16554 ( .A1(n15753), .A2(n15362), .B1(n15795), .B2(n15360), .ZN(
        n15298) );
  AOI211_X1 U16555 ( .C1(n15909), .C2(n15365), .A(n15299), .B(n15298), .ZN(
        n15300) );
  OAI21_X1 U16556 ( .B1(n15301), .B2(n15367), .A(n15300), .ZN(P1_U3228) );
  XOR2_X1 U16557 ( .A(n15303), .B(n15302), .Z(n15308) );
  INV_X1 U16558 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n15304) );
  OAI22_X1 U16559 ( .A1(n15362), .A2(n15579), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15304), .ZN(n15306) );
  OAI22_X1 U16560 ( .A1(n15557), .A2(n15359), .B1(n15360), .B2(n15670), .ZN(
        n15305) );
  AOI211_X1 U16561 ( .C1(n15859), .C2(n15365), .A(n15306), .B(n15305), .ZN(
        n15307) );
  OAI21_X1 U16562 ( .B1(n15308), .B2(n15367), .A(n15307), .ZN(P1_U3229) );
  AOI211_X1 U16563 ( .C1(n15311), .C2(n15310), .A(n15367), .B(n15309), .ZN(
        n15317) );
  INV_X1 U16564 ( .A(n15889), .ZN(n15528) );
  AOI22_X1 U16565 ( .A1(n15337), .A2(n15769), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15315) );
  INV_X1 U16566 ( .A(n15362), .ZN(n15313) );
  AOI22_X1 U16567 ( .A1(n15736), .A2(n15313), .B1(n15740), .B2(n15312), .ZN(
        n15314) );
  OAI211_X1 U16568 ( .C1(n15528), .C2(n15340), .A(n15315), .B(n15314), .ZN(
        n15316) );
  OR2_X1 U16569 ( .A1(n15317), .A2(n15316), .ZN(P1_U3233) );
  INV_X1 U16570 ( .A(n15318), .ZN(n15323) );
  AOI21_X1 U16571 ( .B1(n15320), .B2(n15322), .A(n15319), .ZN(n15321) );
  AOI21_X1 U16572 ( .B1(n15323), .B2(n15322), .A(n15321), .ZN(n15328) );
  INV_X1 U16573 ( .A(n15736), .ZN(n15573) );
  INV_X1 U16574 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n15324) );
  OAI22_X1 U16575 ( .A1(n15573), .A2(n15359), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15324), .ZN(n15326) );
  OAI22_X1 U16576 ( .A1(n15557), .A2(n15362), .B1(n15705), .B2(n15360), .ZN(
        n15325) );
  AOI211_X1 U16577 ( .C1(n15698), .C2(n15365), .A(n15326), .B(n15325), .ZN(
        n15327) );
  OAI21_X1 U16578 ( .B1(n15328), .B2(n15367), .A(n15327), .ZN(P1_U3235) );
  OAI21_X1 U16579 ( .B1(n15331), .B2(n15330), .A(n15329), .ZN(n15333) );
  NAND2_X1 U16580 ( .A1(n15333), .A2(n15332), .ZN(n15339) );
  INV_X1 U16581 ( .A(n15334), .ZN(n15336) );
  INV_X1 U16582 ( .A(n15769), .ZN(n15570) );
  OAI22_X1 U16583 ( .A1(n15570), .A2(n15362), .B1(n15775), .B2(n15360), .ZN(
        n15335) );
  AOI211_X1 U16584 ( .C1(n15337), .C2(n15768), .A(n15336), .B(n15335), .ZN(
        n15338) );
  OAI211_X1 U16585 ( .C1(n15905), .C2(n15340), .A(n15339), .B(n15338), .ZN(
        P1_U3238) );
  INV_X1 U16586 ( .A(n15341), .ZN(n15342) );
  NOR2_X1 U16587 ( .A1(n15343), .A2(n15342), .ZN(n15344) );
  XNOR2_X1 U16588 ( .A(n15345), .B(n15344), .ZN(n15350) );
  INV_X1 U16589 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n15346) );
  OAI22_X1 U16590 ( .A1(n15359), .A2(n15579), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15346), .ZN(n15348) );
  OAI22_X1 U16591 ( .A1(n15362), .A2(n15636), .B1(n15639), .B2(n15360), .ZN(
        n15347) );
  AOI211_X1 U16592 ( .C1(n15847), .C2(n15365), .A(n15348), .B(n15347), .ZN(
        n15349) );
  OAI21_X1 U16593 ( .B1(n15350), .B2(n15367), .A(n15349), .ZN(P1_U3240) );
  INV_X1 U16594 ( .A(n15351), .ZN(n15356) );
  AOI21_X1 U16595 ( .B1(n15353), .B2(n15355), .A(n15352), .ZN(n15354) );
  AOI21_X1 U16596 ( .B1(n15356), .B2(n15355), .A(n15354), .ZN(n15368) );
  OAI21_X1 U16597 ( .B1(n15359), .B2(n15358), .A(n15357), .ZN(n15364) );
  OAI22_X1 U16598 ( .A1(n15362), .A2(n15564), .B1(n15361), .B2(n15360), .ZN(
        n15363) );
  AOI211_X1 U16599 ( .C1(n15561), .C2(n15365), .A(n15364), .B(n15363), .ZN(
        n15366) );
  OAI21_X1 U16600 ( .B1(n15368), .B2(n15367), .A(n15366), .ZN(P1_U3241) );
  MUX2_X1 U16601 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n15531), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16602 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n15586), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16603 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n15369), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16604 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n15613), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16605 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n15370), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16606 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n15614), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16607 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n15667), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16608 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n15577), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16609 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n15703), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16610 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n15554), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16611 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n15736), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16612 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n15550), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16613 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n15769), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16614 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15790), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16615 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n15768), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16616 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n15788), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16617 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n15540), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16618 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n15371), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16619 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n15372), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16620 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n15373), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16621 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n15374), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16622 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n15375), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16623 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n15376), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16624 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n15377), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16625 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n15378), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16626 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n15379), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16627 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n15380), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16628 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n15381), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16629 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n15382), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16630 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n15383), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16631 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n15384), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16632 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n15385), .S(P1_U4016), .Z(
        P1_U3560) );
  AOI211_X1 U16633 ( .C1(n15388), .C2(n15387), .A(n15386), .B(n15398), .ZN(
        n15389) );
  INV_X1 U16634 ( .A(n15389), .ZN(n15397) );
  AOI22_X1 U16635 ( .A1(n16162), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n15396) );
  NAND2_X1 U16636 ( .A1(n15477), .A2(n15390), .ZN(n15395) );
  OAI211_X1 U16637 ( .C1(n15393), .C2(n15392), .A(n15516), .B(n15391), .ZN(
        n15394) );
  NAND4_X1 U16638 ( .A1(n15397), .A2(n15396), .A3(n15395), .A4(n15394), .ZN(
        P1_U3244) );
  AOI22_X1 U16639 ( .A1(n16162), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n15408) );
  AOI211_X1 U16640 ( .C1(n15400), .C2(n15399), .A(n15418), .B(n15398), .ZN(
        n15406) );
  XNOR2_X1 U16641 ( .A(n15402), .B(n15401), .ZN(n15403) );
  OAI22_X1 U16642 ( .A1(n15404), .A2(n15511), .B1(n15512), .B2(n15403), .ZN(
        n15405) );
  NOR2_X1 U16643 ( .A1(n15406), .A2(n15405), .ZN(n15407) );
  NAND3_X1 U16644 ( .A1(n15409), .A2(n15408), .A3(n15407), .ZN(P1_U3245) );
  OAI22_X1 U16645 ( .A1(n15524), .A2(n16192), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15410), .ZN(n15411) );
  AOI21_X1 U16646 ( .B1(n15412), .B2(n15477), .A(n15411), .ZN(n15423) );
  OAI211_X1 U16647 ( .C1(n15415), .C2(n15414), .A(n15516), .B(n15413), .ZN(
        n15422) );
  OR3_X1 U16648 ( .A1(n15418), .A2(n15417), .A3(n15416), .ZN(n15419) );
  NAND3_X1 U16649 ( .A1(n15517), .A2(n15420), .A3(n15419), .ZN(n15421) );
  NAND3_X1 U16650 ( .A1(n15423), .A2(n15422), .A3(n15421), .ZN(P1_U3246) );
  INV_X1 U16651 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n15425) );
  OAI21_X1 U16652 ( .B1(n15524), .B2(n15425), .A(n15424), .ZN(n15426) );
  AOI21_X1 U16653 ( .B1(n15431), .B2(n15477), .A(n15426), .ZN(n15439) );
  OAI21_X1 U16654 ( .B1(n15429), .B2(n15428), .A(n15427), .ZN(n15430) );
  NAND2_X1 U16655 ( .A1(n15517), .A2(n15430), .ZN(n15438) );
  MUX2_X1 U16656 ( .A(n10769), .B(P1_REG2_REG_5__SCAN_IN), .S(n15431), .Z(
        n15432) );
  NAND3_X1 U16657 ( .A1(n15434), .A2(n15433), .A3(n15432), .ZN(n15435) );
  NAND3_X1 U16658 ( .A1(n15516), .A2(n15436), .A3(n15435), .ZN(n15437) );
  NAND3_X1 U16659 ( .A1(n15439), .A2(n15438), .A3(n15437), .ZN(P1_U3248) );
  INV_X1 U16660 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n15441) );
  OAI21_X1 U16661 ( .B1(n15524), .B2(n15441), .A(n15440), .ZN(n15442) );
  AOI21_X1 U16662 ( .B1(n15443), .B2(n15477), .A(n15442), .ZN(n15456) );
  MUX2_X1 U16663 ( .A(n11331), .B(P1_REG2_REG_7__SCAN_IN), .S(n15443), .Z(
        n15444) );
  NAND3_X1 U16664 ( .A1(n15446), .A2(n15445), .A3(n15444), .ZN(n15447) );
  NAND3_X1 U16665 ( .A1(n15516), .A2(n15465), .A3(n15447), .ZN(n15455) );
  INV_X1 U16666 ( .A(n15448), .ZN(n15453) );
  NAND3_X1 U16667 ( .A1(n15451), .A2(n15450), .A3(n15449), .ZN(n15452) );
  NAND3_X1 U16668 ( .A1(n15453), .A2(n15517), .A3(n15452), .ZN(n15454) );
  NAND3_X1 U16669 ( .A1(n15456), .A2(n15455), .A3(n15454), .ZN(P1_U3250) );
  OAI21_X1 U16670 ( .B1(n15458), .B2(n15457), .A(n15472), .ZN(n15459) );
  NAND2_X1 U16671 ( .A1(n15459), .A2(n15517), .ZN(n15469) );
  INV_X1 U16672 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n16234) );
  OAI21_X1 U16673 ( .B1(n15524), .B2(n16234), .A(n15460), .ZN(n15461) );
  AOI21_X1 U16674 ( .B1(n15462), .B2(n15477), .A(n15461), .ZN(n15468) );
  MUX2_X1 U16675 ( .A(n11069), .B(P1_REG2_REG_8__SCAN_IN), .S(n15462), .Z(
        n15463) );
  NAND3_X1 U16676 ( .A1(n15465), .A2(n15464), .A3(n15463), .ZN(n15466) );
  NAND3_X1 U16677 ( .A1(n15516), .A2(n15481), .A3(n15466), .ZN(n15467) );
  NAND3_X1 U16678 ( .A1(n15469), .A2(n15468), .A3(n15467), .ZN(P1_U3251) );
  AND3_X1 U16679 ( .A1(n15472), .A2(n15471), .A3(n15470), .ZN(n15473) );
  OAI21_X1 U16680 ( .B1(n15474), .B2(n15473), .A(n15517), .ZN(n15485) );
  INV_X1 U16681 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n16251) );
  OAI21_X1 U16682 ( .B1(n15524), .B2(n16251), .A(n15475), .ZN(n15476) );
  AOI21_X1 U16683 ( .B1(n15478), .B2(n15477), .A(n15476), .ZN(n15484) );
  MUX2_X1 U16684 ( .A(n11303), .B(P1_REG2_REG_9__SCAN_IN), .S(n15478), .Z(
        n15479) );
  NAND3_X1 U16685 ( .A1(n15481), .A2(n15480), .A3(n15479), .ZN(n15482) );
  NAND3_X1 U16686 ( .A1(n15516), .A2(n15495), .A3(n15482), .ZN(n15483) );
  NAND3_X1 U16687 ( .A1(n15485), .A2(n15484), .A3(n15483), .ZN(P1_U3252) );
  OAI211_X1 U16688 ( .C1(n15488), .C2(n15487), .A(n15486), .B(n15517), .ZN(
        n15500) );
  NOR2_X1 U16689 ( .A1(n15511), .A2(n15489), .ZN(n15490) );
  AOI211_X1 U16690 ( .C1(n16162), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n15491), 
        .B(n15490), .ZN(n15499) );
  MUX2_X1 U16691 ( .A(n11595), .B(P1_REG2_REG_10__SCAN_IN), .S(n15492), .Z(
        n15493) );
  NAND3_X1 U16692 ( .A1(n15495), .A2(n15494), .A3(n15493), .ZN(n15496) );
  NAND3_X1 U16693 ( .A1(n15516), .A2(n15497), .A3(n15496), .ZN(n15498) );
  NAND3_X1 U16694 ( .A1(n15500), .A2(n15499), .A3(n15498), .ZN(P1_U3253) );
  NAND2_X1 U16695 ( .A1(n15507), .A2(n15501), .ZN(n15503) );
  NAND2_X1 U16696 ( .A1(n15503), .A2(n15502), .ZN(n15504) );
  XNOR2_X1 U16697 ( .A(n15505), .B(n15504), .ZN(n15518) );
  INV_X1 U16698 ( .A(n15518), .ZN(n15514) );
  NAND2_X1 U16699 ( .A1(n15507), .A2(n15506), .ZN(n15509) );
  NAND2_X1 U16700 ( .A1(n15509), .A2(n15508), .ZN(n15510) );
  XOR2_X1 U16701 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n15510), .Z(n15515) );
  OAI21_X1 U16702 ( .B1(n15515), .B2(n15512), .A(n15511), .ZN(n15513) );
  AOI21_X1 U16703 ( .B1(n15514), .B2(n15517), .A(n15513), .ZN(n15521) );
  AOI22_X1 U16704 ( .A1(n15518), .A2(n15517), .B1(n15516), .B2(n15515), .ZN(
        n15520) );
  MUX2_X1 U16705 ( .A(n15521), .B(n15520), .S(n15519), .Z(n15523) );
  OAI211_X1 U16706 ( .C1(n15525), .C2(n15524), .A(n15523), .B(n15522), .ZN(
        P1_U3262) );
  NAND2_X1 U16707 ( .A1(n15528), .A2(n15527), .ZN(n15731) );
  OR2_X2 U16708 ( .A1(n15731), .A2(n15883), .ZN(n15718) );
  INV_X1 U16709 ( .A(n15584), .ZN(n15536) );
  NAND2_X1 U16710 ( .A1(n15826), .A2(n15536), .ZN(n15535) );
  XNOR2_X1 U16711 ( .A(n15823), .B(n15535), .ZN(n15529) );
  NAND2_X1 U16712 ( .A1(n15529), .A2(n15910), .ZN(n15822) );
  NOR2_X1 U16713 ( .A1(n15812), .A2(n15530), .ZN(n15532) );
  AOI21_X1 U16714 ( .B1(n16159), .B2(P1_B_REG_SCAN_IN), .A(n16389), .ZN(n15587) );
  NAND2_X1 U16715 ( .A1(n15587), .A2(n15531), .ZN(n15824) );
  NOR2_X1 U16716 ( .A1(n16605), .A2(n15824), .ZN(n15538) );
  AOI211_X1 U16717 ( .C1(n15533), .C2(n16525), .A(n15532), .B(n15538), .ZN(
        n15534) );
  OAI21_X1 U16718 ( .B1(n15822), .B2(n15780), .A(n15534), .ZN(P1_U3263) );
  OAI211_X1 U16719 ( .C1(n15826), .C2(n15536), .A(n15535), .B(n15910), .ZN(
        n15825) );
  NOR2_X1 U16720 ( .A1(n15826), .A2(n16595), .ZN(n15537) );
  AOI211_X1 U16721 ( .C1(n16605), .C2(P1_REG2_REG_30__SCAN_IN), .A(n15538), 
        .B(n15537), .ZN(n15539) );
  OAI21_X1 U16722 ( .B1(n15780), .B2(n15825), .A(n15539), .ZN(P1_U3264) );
  OR2_X1 U16723 ( .A1(n15919), .A2(n15788), .ZN(n15543) );
  NAND2_X1 U16724 ( .A1(n15909), .A2(n15768), .ZN(n15544) );
  NAND2_X1 U16725 ( .A1(n15905), .A2(n15753), .ZN(n15545) );
  NAND2_X1 U16726 ( .A1(n15546), .A2(n15545), .ZN(n15756) );
  OR2_X1 U16727 ( .A1(n15746), .A2(n15769), .ZN(n15548) );
  NAND2_X1 U16728 ( .A1(n15889), .A2(n15550), .ZN(n15551) );
  OR2_X1 U16729 ( .A1(n15883), .A2(n15736), .ZN(n15553) );
  NAND2_X1 U16730 ( .A1(n15724), .A2(n15553), .ZN(n15694) );
  OR2_X1 U16731 ( .A1(n15698), .A2(n15554), .ZN(n15555) );
  INV_X1 U16732 ( .A(n15650), .ZN(n15648) );
  INV_X1 U16733 ( .A(n15847), .ZN(n15580) );
  NAND2_X1 U16734 ( .A1(n15602), .A2(n7811), .ZN(n15601) );
  NAND2_X1 U16735 ( .A1(n15560), .A2(n15559), .ZN(n15563) );
  OR2_X1 U16736 ( .A1(n15561), .A2(n15806), .ZN(n15562) );
  NAND2_X1 U16737 ( .A1(n15563), .A2(n15562), .ZN(n15801) );
  OR2_X2 U16738 ( .A1(n15801), .A2(n15816), .ZN(n15799) );
  NAND2_X1 U16739 ( .A1(n15919), .A2(n15564), .ZN(n15565) );
  NAND2_X1 U16740 ( .A1(n15799), .A2(n15565), .ZN(n15786) );
  OR2_X1 U16741 ( .A1(n15909), .A2(n15807), .ZN(n15566) );
  NAND2_X1 U16742 ( .A1(n15786), .A2(n15566), .ZN(n15568) );
  NAND2_X1 U16743 ( .A1(n15909), .A2(n15807), .ZN(n15567) );
  NAND2_X1 U16744 ( .A1(n15746), .A2(n15570), .ZN(n15571) );
  OR2_X1 U16745 ( .A1(n15889), .A2(n15754), .ZN(n15572) );
  NAND2_X1 U16746 ( .A1(n15735), .A2(n15572), .ZN(n15713) );
  OR2_X1 U16747 ( .A1(n15883), .A2(n15573), .ZN(n15574) );
  INV_X1 U16748 ( .A(n15664), .ZN(n15676) );
  OAI21_X1 U16749 ( .B1(n15581), .B2(n15837), .A(n15596), .ZN(n15583) );
  OAI211_X1 U16750 ( .C1(n15830), .C2(n15585), .A(n15910), .B(n15584), .ZN(
        n15827) );
  NOR2_X1 U16751 ( .A1(n15827), .A2(n15780), .ZN(n15594) );
  NAND2_X1 U16752 ( .A1(n15587), .A2(n15586), .ZN(n15829) );
  OAI22_X1 U16753 ( .A1(n15589), .A2(n15829), .B1(n15588), .B2(n16395), .ZN(
        n15591) );
  NAND2_X1 U16754 ( .A1(n15787), .A2(n15613), .ZN(n15828) );
  NOR2_X1 U16755 ( .A1(n16605), .A2(n15828), .ZN(n15590) );
  AOI211_X1 U16756 ( .C1(n16605), .C2(P1_REG2_REG_29__SCAN_IN), .A(n15591), 
        .B(n15590), .ZN(n15592) );
  OAI21_X1 U16757 ( .B1(n15830), .B2(n16595), .A(n15592), .ZN(n15593) );
  AOI211_X1 U16758 ( .C1(n15832), .C2(n15711), .A(n15594), .B(n15593), .ZN(
        n15595) );
  OAI21_X1 U16759 ( .B1(n15834), .B2(n16597), .A(n15595), .ZN(P1_U3356) );
  OAI211_X1 U16760 ( .C1(n15598), .C2(n15597), .A(n15596), .B(n16458), .ZN(
        n15600) );
  OAI21_X1 U16761 ( .B1(n15602), .B2(n7811), .A(n15601), .ZN(n15838) );
  INV_X1 U16762 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n15604) );
  OAI22_X1 U16763 ( .A1(n15812), .A2(n15604), .B1(n15603), .B2(n16395), .ZN(
        n15605) );
  AOI21_X1 U16764 ( .B1(n15837), .B2(n16525), .A(n15605), .ZN(n15609) );
  NAND2_X1 U16765 ( .A1(n15837), .A2(n15615), .ZN(n15606) );
  NAND2_X1 U16766 ( .A1(n15836), .A2(n16601), .ZN(n15608) );
  OAI211_X1 U16767 ( .C1(n15838), .C2(n16597), .A(n15609), .B(n15608), .ZN(
        n15610) );
  AOI21_X1 U16768 ( .B1(n15835), .B2(n15812), .A(n15610), .ZN(n15611) );
  INV_X1 U16769 ( .A(n15611), .ZN(P1_U3265) );
  INV_X1 U16770 ( .A(n15635), .ZN(n15617) );
  INV_X1 U16771 ( .A(n15615), .ZN(n15616) );
  AOI211_X1 U16772 ( .C1(n15840), .C2(n15617), .A(n15915), .B(n15616), .ZN(
        n15839) );
  INV_X1 U16773 ( .A(n15618), .ZN(n15619) );
  AOI22_X1 U16774 ( .A1(n16605), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n15619), 
        .B2(n16592), .ZN(n15620) );
  OAI21_X1 U16775 ( .B1(n15621), .B2(n16595), .A(n15620), .ZN(n15626) );
  AOI21_X1 U16776 ( .B1(n15624), .B2(n15623), .A(n15622), .ZN(n15843) );
  NOR2_X1 U16777 ( .A1(n15843), .A2(n16597), .ZN(n15625) );
  AOI211_X1 U16778 ( .C1(n15839), .C2(n16601), .A(n15626), .B(n15625), .ZN(
        n15627) );
  OAI21_X1 U16779 ( .B1(n15842), .B2(n16605), .A(n15627), .ZN(P1_U3266) );
  OAI21_X1 U16780 ( .B1(n15629), .B2(n15630), .A(n15628), .ZN(n15850) );
  XNOR2_X1 U16781 ( .A(n15631), .B(n15630), .ZN(n15844) );
  NAND2_X1 U16782 ( .A1(n15844), .A2(n15711), .ZN(n15646) );
  NAND2_X1 U16783 ( .A1(n15847), .A2(n15632), .ZN(n15633) );
  NAND2_X1 U16784 ( .A1(n15633), .A2(n15910), .ZN(n15634) );
  NOR2_X1 U16785 ( .A1(n15635), .A2(n15634), .ZN(n15845) );
  NAND2_X1 U16786 ( .A1(n15847), .A2(n16525), .ZN(n15642) );
  OR2_X1 U16787 ( .A1(n15636), .A2(n16389), .ZN(n15638) );
  NAND2_X1 U16788 ( .A1(n15787), .A2(n15667), .ZN(n15637) );
  NAND2_X1 U16789 ( .A1(n15638), .A2(n15637), .ZN(n15846) );
  NOR2_X1 U16790 ( .A1(n16395), .A2(n15639), .ZN(n15640) );
  AOI21_X1 U16791 ( .B1(n15812), .B2(n15846), .A(n15640), .ZN(n15641) );
  OAI211_X1 U16792 ( .C1(n15812), .C2(n15643), .A(n15642), .B(n15641), .ZN(
        n15644) );
  AOI21_X1 U16793 ( .B1(n15845), .B2(n16601), .A(n15644), .ZN(n15645) );
  OAI211_X1 U16794 ( .C1(n15850), .C2(n16597), .A(n15646), .B(n15645), .ZN(
        P1_U3267) );
  OAI21_X1 U16795 ( .B1(n15649), .B2(n15648), .A(n15647), .ZN(n15856) );
  XNOR2_X1 U16796 ( .A(n15651), .B(n15650), .ZN(n15851) );
  NAND2_X1 U16797 ( .A1(n15851), .A2(n15711), .ZN(n15661) );
  XNOR2_X1 U16798 ( .A(n15853), .B(n15665), .ZN(n15654) );
  OAI222_X1 U16799 ( .A1(n15654), .A2(n15915), .B1(n16389), .B2(n15653), .C1(
        n15805), .C2(n15652), .ZN(n15852) );
  NOR2_X1 U16800 ( .A1(n15655), .A2(n16595), .ZN(n15659) );
  INV_X1 U16801 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n15657) );
  OAI22_X1 U16802 ( .A1(n15812), .A2(n15657), .B1(n15656), .B2(n16395), .ZN(
        n15658) );
  AOI211_X1 U16803 ( .C1(n15852), .C2(n16601), .A(n15659), .B(n15658), .ZN(
        n15660) );
  OAI211_X1 U16804 ( .C1(n15856), .C2(n16597), .A(n15661), .B(n15660), .ZN(
        P1_U3268) );
  AOI21_X1 U16805 ( .B1(n15664), .B2(n15663), .A(n15662), .ZN(n15864) );
  AOI21_X1 U16806 ( .B1(n15685), .B2(n15859), .A(n15915), .ZN(n15666) );
  AND2_X1 U16807 ( .A1(n15666), .A2(n15665), .ZN(n15857) );
  NAND2_X1 U16808 ( .A1(n15859), .A2(n16525), .ZN(n15674) );
  NAND2_X1 U16809 ( .A1(n15703), .A2(n15787), .ZN(n15669) );
  NAND2_X1 U16810 ( .A1(n15789), .A2(n15667), .ZN(n15668) );
  NAND2_X1 U16811 ( .A1(n15669), .A2(n15668), .ZN(n15858) );
  INV_X1 U16812 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n15671) );
  OAI22_X1 U16813 ( .A1(n15812), .A2(n15671), .B1(n15670), .B2(n16395), .ZN(
        n15672) );
  AOI21_X1 U16814 ( .B1(n15858), .B2(n15812), .A(n15672), .ZN(n15673) );
  NAND2_X1 U16815 ( .A1(n15674), .A2(n15673), .ZN(n15675) );
  AOI21_X1 U16816 ( .B1(n15857), .B2(n16601), .A(n15675), .ZN(n15679) );
  NAND2_X1 U16817 ( .A1(n15677), .A2(n15676), .ZN(n15860) );
  NAND3_X1 U16818 ( .A1(n15861), .A2(n15711), .A3(n15860), .ZN(n15678) );
  OAI211_X1 U16819 ( .C1(n15864), .C2(n16597), .A(n15679), .B(n15678), .ZN(
        P1_U3269) );
  XNOR2_X1 U16820 ( .A(n15680), .B(n15556), .ZN(n15681) );
  NAND2_X1 U16821 ( .A1(n15681), .A2(n16458), .ZN(n15683) );
  NAND2_X1 U16822 ( .A1(n15683), .A2(n15682), .ZN(n15872) );
  AOI21_X1 U16823 ( .B1(n15684), .B2(n16592), .A(n15872), .ZN(n15693) );
  OAI211_X1 U16824 ( .C1(n15686), .C2(n15701), .A(n15910), .B(n15685), .ZN(
        n15869) );
  NAND2_X1 U16825 ( .A1(n15688), .A2(n15687), .ZN(n15865) );
  NAND3_X1 U16826 ( .A1(n15866), .A2(n15865), .A3(n15818), .ZN(n15690) );
  AOI22_X1 U16827 ( .A1(n15867), .A2(n16525), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n16605), .ZN(n15689) );
  OAI211_X1 U16828 ( .C1(n15869), .C2(n15780), .A(n15690), .B(n15689), .ZN(
        n15691) );
  INV_X1 U16829 ( .A(n15691), .ZN(n15692) );
  OAI21_X1 U16830 ( .B1(n15693), .B2(n16605), .A(n15692), .ZN(P1_U3270) );
  XNOR2_X1 U16831 ( .A(n15694), .B(n15696), .ZN(n15881) );
  OAI21_X1 U16832 ( .B1(n15697), .B2(n15696), .A(n15695), .ZN(n15879) );
  NAND2_X1 U16833 ( .A1(n15698), .A2(n15718), .ZN(n15699) );
  NAND2_X1 U16834 ( .A1(n15699), .A2(n15910), .ZN(n15700) );
  NOR2_X1 U16835 ( .A1(n15701), .A2(n15700), .ZN(n15878) );
  NAND2_X1 U16836 ( .A1(n15878), .A2(n16601), .ZN(n15709) );
  AND2_X1 U16837 ( .A1(n15736), .A2(n15787), .ZN(n15702) );
  AOI21_X1 U16838 ( .B1(n15703), .B2(n15789), .A(n15702), .ZN(n15875) );
  INV_X1 U16839 ( .A(n15875), .ZN(n15707) );
  INV_X1 U16840 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n15704) );
  OAI22_X1 U16841 ( .A1(n15705), .A2(n16395), .B1(n15704), .B2(n15812), .ZN(
        n15706) );
  AOI21_X1 U16842 ( .B1(n15707), .B2(n15812), .A(n15706), .ZN(n15708) );
  OAI211_X1 U16843 ( .C1(n16595), .C2(n15876), .A(n15709), .B(n15708), .ZN(
        n15710) );
  AOI21_X1 U16844 ( .B1(n15879), .B2(n15711), .A(n15710), .ZN(n15712) );
  OAI21_X1 U16845 ( .B1(n15881), .B2(n16597), .A(n15712), .ZN(P1_U3271) );
  INV_X1 U16846 ( .A(n15713), .ZN(n15714) );
  AOI21_X1 U16847 ( .B1(n15714), .B2(n7873), .A(n16558), .ZN(n15717) );
  AOI21_X1 U16848 ( .B1(n15717), .B2(n15716), .A(n15715), .ZN(n15885) );
  INV_X1 U16849 ( .A(n15718), .ZN(n15719) );
  AOI211_X1 U16850 ( .C1(n15883), .C2(n15731), .A(n15915), .B(n15719), .ZN(
        n15882) );
  INV_X1 U16851 ( .A(n15720), .ZN(n15721) );
  AOI22_X1 U16852 ( .A1(n15721), .A2(n16592), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n16605), .ZN(n15722) );
  OAI21_X1 U16853 ( .B1(n15723), .B2(n16595), .A(n15722), .ZN(n15728) );
  AOI21_X1 U16854 ( .B1(n15726), .B2(n15725), .A(n15552), .ZN(n15886) );
  NOR2_X1 U16855 ( .A1(n15886), .A2(n16597), .ZN(n15727) );
  AOI211_X1 U16856 ( .C1(n15882), .C2(n16601), .A(n15728), .B(n15727), .ZN(
        n15729) );
  OAI21_X1 U16857 ( .B1(n16605), .B2(n15885), .A(n15729), .ZN(P1_U3272) );
  NAND2_X1 U16858 ( .A1(n15889), .A2(n15748), .ZN(n15730) );
  AND2_X1 U16859 ( .A1(n15731), .A2(n15730), .ZN(n15890) );
  INV_X1 U16860 ( .A(n15890), .ZN(n15732) );
  NOR2_X1 U16861 ( .A1(n15732), .A2(n15810), .ZN(n15739) );
  NAND2_X1 U16862 ( .A1(n15733), .A2(n15549), .ZN(n15734) );
  NAND3_X1 U16863 ( .A1(n15735), .A2(n16458), .A3(n15734), .ZN(n15738) );
  AOI22_X1 U16864 ( .A1(n15736), .A2(n15789), .B1(n15787), .B2(n15769), .ZN(
        n15737) );
  NAND2_X1 U16865 ( .A1(n15738), .A2(n15737), .ZN(n15894) );
  AOI211_X1 U16866 ( .C1(n16592), .C2(n15740), .A(n15739), .B(n15894), .ZN(
        n15745) );
  AOI22_X1 U16867 ( .A1(n15889), .A2(n16525), .B1(n16605), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n15744) );
  NAND2_X1 U16868 ( .A1(n15742), .A2(n15741), .ZN(n15887) );
  NAND3_X1 U16869 ( .A1(n15888), .A2(n15887), .A3(n15818), .ZN(n15743) );
  OAI211_X1 U16870 ( .C1(n15745), .C2(n16605), .A(n15744), .B(n15743), .ZN(
        P1_U3273) );
  INV_X1 U16871 ( .A(n15810), .ZN(n15793) );
  NAND2_X1 U16872 ( .A1(n15774), .A2(n15746), .ZN(n15747) );
  NAND2_X1 U16873 ( .A1(n15748), .A2(n15747), .ZN(n15898) );
  INV_X1 U16874 ( .A(n15898), .ZN(n15755) );
  INV_X1 U16875 ( .A(n15749), .ZN(n15750) );
  AOI21_X1 U16876 ( .B1(n15757), .B2(n15751), .A(n15750), .ZN(n15752) );
  OAI222_X1 U16877 ( .A1(n16389), .A2(n15754), .B1(n15805), .B2(n15753), .C1(
        n16558), .C2(n15752), .ZN(n15899) );
  AOI21_X1 U16878 ( .B1(n15793), .B2(n15755), .A(n15899), .ZN(n15762) );
  XNOR2_X1 U16879 ( .A(n15756), .B(n15757), .ZN(n15901) );
  AOI22_X1 U16880 ( .A1(n16605), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n15758), 
        .B2(n16592), .ZN(n15759) );
  OAI21_X1 U16881 ( .B1(n15897), .B2(n16595), .A(n15759), .ZN(n15760) );
  AOI21_X1 U16882 ( .B1(n15901), .B2(n15818), .A(n15760), .ZN(n15761) );
  OAI21_X1 U16883 ( .B1(n15762), .B2(n16605), .A(n15761), .ZN(P1_U3274) );
  XNOR2_X1 U16884 ( .A(n15763), .B(n15764), .ZN(n15903) );
  INV_X1 U16885 ( .A(n15903), .ZN(n15783) );
  NAND2_X1 U16886 ( .A1(n15765), .A2(n15764), .ZN(n15766) );
  NAND3_X1 U16887 ( .A1(n15767), .A2(n16458), .A3(n15766), .ZN(n15771) );
  AOI22_X1 U16888 ( .A1(n15769), .A2(n15789), .B1(n15787), .B2(n15768), .ZN(
        n15770) );
  NAND2_X1 U16889 ( .A1(n15771), .A2(n15770), .ZN(n15907) );
  INV_X1 U16890 ( .A(n15792), .ZN(n15772) );
  AOI21_X1 U16891 ( .B1(n15778), .B2(n15772), .A(n15915), .ZN(n15773) );
  NAND2_X1 U16892 ( .A1(n15774), .A2(n15773), .ZN(n15904) );
  OAI22_X1 U16893 ( .A1(n15812), .A2(n15776), .B1(n15775), .B2(n16395), .ZN(
        n15777) );
  AOI21_X1 U16894 ( .B1(n15778), .B2(n16525), .A(n15777), .ZN(n15779) );
  OAI21_X1 U16895 ( .B1(n15904), .B2(n15780), .A(n15779), .ZN(n15781) );
  AOI21_X1 U16896 ( .B1(n15907), .B2(n15812), .A(n15781), .ZN(n15782) );
  OAI21_X1 U16897 ( .B1(n16597), .B2(n15783), .A(n15782), .ZN(P1_U3275) );
  XOR2_X1 U16898 ( .A(n15784), .B(n15785), .Z(n15914) );
  XOR2_X1 U16899 ( .A(n15786), .B(n15785), .Z(n15791) );
  AOI222_X1 U16900 ( .A1(n16458), .A2(n15791), .B1(n15790), .B2(n15789), .C1(
        n15788), .C2(n15787), .ZN(n15913) );
  AOI21_X1 U16901 ( .B1(n15909), .B2(n15803), .A(n15792), .ZN(n15911) );
  NAND2_X1 U16902 ( .A1(n15911), .A2(n15793), .ZN(n15794) );
  OAI211_X1 U16903 ( .C1(n16395), .C2(n15795), .A(n15913), .B(n15794), .ZN(
        n15796) );
  NAND2_X1 U16904 ( .A1(n15796), .A2(n15812), .ZN(n15798) );
  AOI22_X1 U16905 ( .A1(n15909), .A2(n16525), .B1(P1_REG2_REG_17__SCAN_IN), 
        .B2(n16605), .ZN(n15797) );
  OAI211_X1 U16906 ( .C1(n15914), .C2(n16597), .A(n15798), .B(n15797), .ZN(
        P1_U3276) );
  INV_X1 U16907 ( .A(n15799), .ZN(n15800) );
  AOI21_X1 U16908 ( .B1(n15816), .B2(n15801), .A(n15800), .ZN(n15923) );
  OAI21_X1 U16909 ( .B1(n7596), .B2(n7597), .A(n15803), .ZN(n15916) );
  INV_X1 U16910 ( .A(n15804), .ZN(n15808) );
  OAI22_X1 U16911 ( .A1(n15807), .A2(n16389), .B1(n15806), .B2(n15805), .ZN(
        n15918) );
  AOI21_X1 U16912 ( .B1(n15808), .B2(n16592), .A(n15918), .ZN(n15809) );
  OAI21_X1 U16913 ( .B1(n15916), .B2(n15810), .A(n15809), .ZN(n15814) );
  INV_X1 U16914 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n15811) );
  OAI22_X1 U16915 ( .A1(n7596), .A2(n16595), .B1(n15812), .B2(n15811), .ZN(
        n15813) );
  AOI21_X1 U16916 ( .B1(n15814), .B2(n15812), .A(n15813), .ZN(n15820) );
  OAI21_X1 U16917 ( .B1(n15817), .B2(n15816), .A(n15815), .ZN(n15920) );
  NAND2_X1 U16918 ( .A1(n15920), .A2(n15818), .ZN(n15819) );
  OAI211_X1 U16919 ( .C1(n15923), .C2(n15821), .A(n15820), .B(n15819), .ZN(
        P1_U3277) );
  OAI211_X1 U16920 ( .C1(n15823), .C2(n16556), .A(n15822), .B(n15824), .ZN(
        n15946) );
  MUX2_X1 U16921 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15946), .S(n16469), .Z(
        P1_U3559) );
  OAI211_X1 U16922 ( .C1(n15826), .C2(n16556), .A(n15825), .B(n15824), .ZN(
        n15947) );
  MUX2_X1 U16923 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15947), .S(n16469), .Z(
        P1_U3558) );
  OAI211_X1 U16924 ( .C1(n15830), .C2(n16556), .A(n15829), .B(n15828), .ZN(
        n15831) );
  MUX2_X1 U16925 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15948), .S(n16469), .Z(
        P1_U3556) );
  AOI21_X1 U16926 ( .B1(n16490), .B2(n15840), .A(n15839), .ZN(n15841) );
  MUX2_X1 U16927 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15949), .S(n16469), .Z(
        P1_U3555) );
  NAND2_X1 U16928 ( .A1(n15844), .A2(n16458), .ZN(n15849) );
  AOI211_X1 U16929 ( .C1(n16490), .C2(n15847), .A(n15846), .B(n15845), .ZN(
        n15848) );
  OAI211_X1 U16930 ( .C1(n16435), .C2(n15850), .A(n15849), .B(n15848), .ZN(
        n15950) );
  MUX2_X1 U16931 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15950), .S(n16469), .Z(
        P1_U3554) );
  NAND2_X1 U16932 ( .A1(n15851), .A2(n16458), .ZN(n15855) );
  AOI21_X1 U16933 ( .B1(n16490), .B2(n15853), .A(n15852), .ZN(n15854) );
  OAI211_X1 U16934 ( .C1(n16435), .C2(n15856), .A(n15855), .B(n15854), .ZN(
        n15951) );
  MUX2_X1 U16935 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15951), .S(n16469), .Z(
        P1_U3553) );
  AOI211_X1 U16936 ( .C1(n16490), .C2(n15859), .A(n15858), .B(n15857), .ZN(
        n15863) );
  NAND3_X1 U16937 ( .A1(n15861), .A2(n16458), .A3(n15860), .ZN(n15862) );
  OAI211_X1 U16938 ( .C1(n15864), .C2(n16435), .A(n15863), .B(n15862), .ZN(
        n15952) );
  MUX2_X1 U16939 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15952), .S(n16469), .Z(
        P1_U3552) );
  NAND3_X1 U16940 ( .A1(n15866), .A2(n16564), .A3(n15865), .ZN(n15870) );
  NAND2_X1 U16941 ( .A1(n15867), .A2(n16490), .ZN(n15868) );
  NAND3_X1 U16942 ( .A1(n15870), .A2(n15869), .A3(n15868), .ZN(n15871) );
  NOR2_X1 U16943 ( .A1(n15872), .A2(n15871), .ZN(n15953) );
  MUX2_X1 U16944 ( .A(n15873), .B(n15953), .S(n16469), .Z(n15874) );
  INV_X1 U16945 ( .A(n15874), .ZN(P1_U3551) );
  OAI21_X1 U16946 ( .B1(n15876), .B2(n16556), .A(n15875), .ZN(n15877) );
  AOI211_X1 U16947 ( .C1(n15879), .C2(n16458), .A(n15878), .B(n15877), .ZN(
        n15880) );
  OAI21_X1 U16948 ( .B1(n16435), .B2(n15881), .A(n15880), .ZN(n15956) );
  MUX2_X1 U16949 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15956), .S(n16469), .Z(
        P1_U3550) );
  AOI21_X1 U16950 ( .B1(n16490), .B2(n15883), .A(n15882), .ZN(n15884) );
  OAI211_X1 U16951 ( .C1(n15886), .C2(n16435), .A(n15885), .B(n15884), .ZN(
        n15957) );
  MUX2_X1 U16952 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15957), .S(n16469), .Z(
        P1_U3549) );
  NAND3_X1 U16953 ( .A1(n15888), .A2(n15887), .A3(n16564), .ZN(n15892) );
  AOI22_X1 U16954 ( .A1(n15890), .A2(n15910), .B1(n16490), .B2(n15889), .ZN(
        n15891) );
  NAND2_X1 U16955 ( .A1(n15892), .A2(n15891), .ZN(n15893) );
  NOR2_X1 U16956 ( .A1(n15894), .A2(n15893), .ZN(n15958) );
  MUX2_X1 U16957 ( .A(n15895), .B(n15958), .S(n16469), .Z(n15896) );
  INV_X1 U16958 ( .A(n15896), .ZN(P1_U3548) );
  OAI22_X1 U16959 ( .A1(n15898), .A2(n15915), .B1(n15897), .B2(n16556), .ZN(
        n15900) );
  AOI211_X1 U16960 ( .C1(n15901), .C2(n16564), .A(n15900), .B(n15899), .ZN(
        n15902) );
  INV_X1 U16961 ( .A(n15902), .ZN(n15961) );
  MUX2_X1 U16962 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15961), .S(n16469), .Z(
        P1_U3547) );
  AND2_X1 U16963 ( .A1(n15903), .A2(n16564), .ZN(n15908) );
  OAI21_X1 U16964 ( .B1(n15905), .B2(n16556), .A(n15904), .ZN(n15906) );
  MUX2_X1 U16965 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15962), .S(n16469), .Z(
        P1_U3546) );
  AOI22_X1 U16966 ( .A1(n15911), .A2(n15910), .B1(n16490), .B2(n15909), .ZN(
        n15912) );
  OAI211_X1 U16967 ( .C1(n16435), .C2(n15914), .A(n15913), .B(n15912), .ZN(
        n15963) );
  MUX2_X1 U16968 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15963), .S(n16469), .Z(
        P1_U3545) );
  NOR2_X1 U16969 ( .A1(n15916), .A2(n15915), .ZN(n15917) );
  AOI211_X1 U16970 ( .C1(n16490), .C2(n15919), .A(n15918), .B(n15917), .ZN(
        n15922) );
  NAND2_X1 U16971 ( .A1(n15920), .A2(n16564), .ZN(n15921) );
  OAI211_X1 U16972 ( .C1(n15923), .C2(n16558), .A(n15922), .B(n15921), .ZN(
        n15964) );
  MUX2_X1 U16973 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15964), .S(n16469), .Z(
        P1_U3544) );
  OAI211_X1 U16974 ( .C1(n15926), .C2(n16556), .A(n15925), .B(n15924), .ZN(
        n15927) );
  AOI21_X1 U16975 ( .B1(n15928), .B2(n16458), .A(n15927), .ZN(n15929) );
  OAI21_X1 U16976 ( .B1(n16435), .B2(n15930), .A(n15929), .ZN(n15965) );
  MUX2_X1 U16977 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15965), .S(n16469), .Z(
        P1_U3543) );
  OAI211_X1 U16978 ( .C1(n15933), .C2(n16556), .A(n15932), .B(n15931), .ZN(
        n15934) );
  AOI21_X1 U16979 ( .B1(n15935), .B2(n16564), .A(n15934), .ZN(n15936) );
  OAI21_X1 U16980 ( .B1(n16558), .B2(n15937), .A(n15936), .ZN(n15966) );
  MUX2_X1 U16981 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15966), .S(n16469), .Z(
        P1_U3542) );
  AOI211_X1 U16982 ( .C1(n16490), .C2(n15940), .A(n15939), .B(n15938), .ZN(
        n15943) );
  NAND2_X1 U16983 ( .A1(n15941), .A2(n16564), .ZN(n15942) );
  OAI211_X1 U16984 ( .C1(n15944), .C2(n16558), .A(n15943), .B(n15942), .ZN(
        n15967) );
  MUX2_X1 U16985 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15967), .S(n16469), .Z(
        P1_U3541) );
  MUX2_X1 U16986 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n15945), .S(n16469), .Z(
        P1_U3533) );
  MUX2_X1 U16987 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15946), .S(n16570), .Z(
        P1_U3527) );
  MUX2_X1 U16988 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15947), .S(n16570), .Z(
        P1_U3526) );
  MUX2_X1 U16989 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15950), .S(n16570), .Z(
        P1_U3522) );
  MUX2_X1 U16990 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15951), .S(n16570), .Z(
        P1_U3521) );
  MUX2_X1 U16991 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15952), .S(n16570), .Z(
        P1_U3520) );
  INV_X1 U16992 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n15954) );
  MUX2_X1 U16993 ( .A(n15954), .B(n15953), .S(n16570), .Z(n15955) );
  INV_X1 U16994 ( .A(n15955), .ZN(P1_U3519) );
  MUX2_X1 U16995 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15956), .S(n16570), .Z(
        P1_U3518) );
  MUX2_X1 U16996 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15957), .S(n16570), .Z(
        P1_U3517) );
  INV_X1 U16997 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n15959) );
  MUX2_X1 U16998 ( .A(n15959), .B(n15958), .S(n16570), .Z(n15960) );
  INV_X1 U16999 ( .A(n15960), .ZN(P1_U3516) );
  MUX2_X1 U17000 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15961), .S(n16570), .Z(
        P1_U3515) );
  MUX2_X1 U17001 ( .A(n15962), .B(P1_REG0_REG_18__SCAN_IN), .S(n16567), .Z(
        P1_U3513) );
  MUX2_X1 U17002 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15963), .S(n16570), .Z(
        P1_U3510) );
  MUX2_X1 U17003 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15964), .S(n16570), .Z(
        P1_U3507) );
  MUX2_X1 U17004 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15965), .S(n16570), .Z(
        P1_U3504) );
  MUX2_X1 U17005 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15966), .S(n16570), .Z(
        P1_U3501) );
  MUX2_X1 U17006 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n15967), .S(n16570), .Z(
        P1_U3498) );
  MUX2_X1 U17007 ( .A(n15968), .B(P1_D_REG_1__SCAN_IN), .S(n16000), .Z(
        P1_U3446) );
  NOR4_X1 U17008 ( .A1(n15969), .A2(P1_IR_REG_30__SCAN_IN), .A3(n10344), .A4(
        P1_U3086), .ZN(n15970) );
  AOI21_X1 U17009 ( .B1(n15971), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15970), 
        .ZN(n15972) );
  OAI21_X1 U17010 ( .B1(n15973), .B2(n15990), .A(n15972), .ZN(P1_U3324) );
  OAI222_X1 U17011 ( .A1(P1_U3086), .A2(n15979), .B1(n15990), .B2(n15978), 
        .C1(n15977), .C2(n15992), .ZN(P1_U3326) );
  OAI222_X1 U17012 ( .A1(n15982), .A2(P1_U3086), .B1(n15990), .B2(n15981), 
        .C1(n15980), .C2(n15987), .ZN(P1_U3328) );
  OAI222_X1 U17013 ( .A1(P1_U3086), .A2(n15985), .B1(n15990), .B2(n15984), 
        .C1(n15983), .C2(n15992), .ZN(P1_U3329) );
  OAI222_X1 U17014 ( .A1(n15991), .A2(P1_U3086), .B1(n15990), .B2(n15989), 
        .C1(n15988), .C2(n15987), .ZN(P1_U3330) );
  OAI222_X1 U17015 ( .A1(n15995), .A2(P1_U3086), .B1(n15990), .B2(n15994), 
        .C1(n15993), .C2(n15992), .ZN(P1_U3331) );
  MUX2_X1 U17016 ( .A(n15997), .B(n15996), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U17017 ( .A(n15998), .ZN(n15999) );
  MUX2_X1 U17018 ( .A(n15999), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U17019 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n16001) );
  NOR2_X1 U17020 ( .A1(n16031), .A2(n16001), .ZN(P1_U3323) );
  INV_X1 U17021 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n16002) );
  NOR2_X1 U17022 ( .A1(n16031), .A2(n16002), .ZN(P1_U3322) );
  INV_X1 U17023 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n16003) );
  NOR2_X1 U17024 ( .A1(n16031), .A2(n16003), .ZN(P1_U3321) );
  INV_X1 U17025 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n16004) );
  NOR2_X1 U17026 ( .A1(n16031), .A2(n16004), .ZN(P1_U3320) );
  INV_X1 U17027 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n16005) );
  NOR2_X1 U17028 ( .A1(n16031), .A2(n16005), .ZN(P1_U3319) );
  INV_X1 U17029 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n16006) );
  NOR2_X1 U17030 ( .A1(n16031), .A2(n16006), .ZN(P1_U3318) );
  INV_X1 U17031 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n16007) );
  NOR2_X1 U17032 ( .A1(n16031), .A2(n16007), .ZN(P1_U3317) );
  INV_X1 U17033 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n16008) );
  NOR2_X1 U17034 ( .A1(n16031), .A2(n16008), .ZN(P1_U3316) );
  INV_X1 U17035 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n16009) );
  NOR2_X1 U17036 ( .A1(n16031), .A2(n16009), .ZN(P1_U3315) );
  INV_X1 U17037 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n16010) );
  NOR2_X1 U17038 ( .A1(n16031), .A2(n16010), .ZN(P1_U3314) );
  INV_X1 U17039 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n16011) );
  NOR2_X1 U17040 ( .A1(n16031), .A2(n16011), .ZN(P1_U3313) );
  INV_X1 U17041 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n16012) );
  NOR2_X1 U17042 ( .A1(n16031), .A2(n16012), .ZN(P1_U3312) );
  INV_X1 U17043 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n16013) );
  NOR2_X1 U17044 ( .A1(n16031), .A2(n16013), .ZN(P1_U3311) );
  INV_X1 U17045 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n16014) );
  NOR2_X1 U17046 ( .A1(n16031), .A2(n16014), .ZN(P1_U3310) );
  INV_X1 U17047 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n16015) );
  NOR2_X1 U17048 ( .A1(n16031), .A2(n16015), .ZN(P1_U3309) );
  INV_X1 U17049 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n16016) );
  NOR2_X1 U17050 ( .A1(n16031), .A2(n16016), .ZN(P1_U3308) );
  INV_X1 U17051 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n16017) );
  NOR2_X1 U17052 ( .A1(n16031), .A2(n16017), .ZN(P1_U3307) );
  INV_X1 U17053 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n16018) );
  NOR2_X1 U17054 ( .A1(n16031), .A2(n16018), .ZN(P1_U3306) );
  INV_X1 U17055 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n16019) );
  NOR2_X1 U17056 ( .A1(n16031), .A2(n16019), .ZN(P1_U3305) );
  INV_X1 U17057 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n16020) );
  NOR2_X1 U17058 ( .A1(n16031), .A2(n16020), .ZN(P1_U3304) );
  INV_X1 U17059 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n16021) );
  NOR2_X1 U17060 ( .A1(n16031), .A2(n16021), .ZN(P1_U3303) );
  INV_X1 U17061 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n16022) );
  NOR2_X1 U17062 ( .A1(n16031), .A2(n16022), .ZN(P1_U3302) );
  INV_X1 U17063 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n16023) );
  NOR2_X1 U17064 ( .A1(n16031), .A2(n16023), .ZN(P1_U3301) );
  INV_X1 U17065 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n16024) );
  NOR2_X1 U17066 ( .A1(n16031), .A2(n16024), .ZN(P1_U3300) );
  INV_X1 U17067 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n16025) );
  NOR2_X1 U17068 ( .A1(n16031), .A2(n16025), .ZN(P1_U3299) );
  INV_X1 U17069 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n16026) );
  NOR2_X1 U17070 ( .A1(n16031), .A2(n16026), .ZN(P1_U3298) );
  INV_X1 U17071 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n16027) );
  NOR2_X1 U17072 ( .A1(n16031), .A2(n16027), .ZN(P1_U3297) );
  INV_X1 U17073 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n16028) );
  NOR2_X1 U17074 ( .A1(n16031), .A2(n16028), .ZN(P1_U3296) );
  INV_X1 U17075 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n16029) );
  NOR2_X1 U17076 ( .A1(n16031), .A2(n16029), .ZN(P1_U3295) );
  INV_X1 U17077 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n16030) );
  NOR2_X1 U17078 ( .A1(n16031), .A2(n16030), .ZN(P1_U3294) );
  INV_X1 U17079 ( .A(n16040), .ZN(n16037) );
  AOI21_X1 U17080 ( .B1(n16033), .B2(n16037), .A(n16032), .ZN(P2_U3417) );
  AND2_X1 U17081 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n16035), .ZN(P2_U3295) );
  AND2_X1 U17082 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n16035), .ZN(P2_U3294) );
  AND2_X1 U17083 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n16035), .ZN(P2_U3293) );
  AND2_X1 U17084 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n16035), .ZN(P2_U3292) );
  AND2_X1 U17085 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n16035), .ZN(P2_U3291) );
  AND2_X1 U17086 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n16035), .ZN(P2_U3290) );
  AND2_X1 U17087 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n16035), .ZN(P2_U3289) );
  AND2_X1 U17088 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n16035), .ZN(P2_U3288) );
  AND2_X1 U17089 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n16035), .ZN(P2_U3287) );
  AND2_X1 U17090 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n16035), .ZN(P2_U3286) );
  AND2_X1 U17091 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n16035), .ZN(P2_U3285) );
  AND2_X1 U17092 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n16035), .ZN(P2_U3284) );
  AND2_X1 U17093 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n16035), .ZN(P2_U3283) );
  AND2_X1 U17094 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n16035), .ZN(P2_U3282) );
  AND2_X1 U17095 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n16035), .ZN(P2_U3281) );
  AND2_X1 U17096 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n16035), .ZN(P2_U3280) );
  AND2_X1 U17097 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n16035), .ZN(P2_U3279) );
  AND2_X1 U17098 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n16035), .ZN(P2_U3278) );
  AND2_X1 U17099 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n16035), .ZN(P2_U3277) );
  AND2_X1 U17100 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n16035), .ZN(P2_U3276) );
  AND2_X1 U17101 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n16035), .ZN(P2_U3275) );
  AND2_X1 U17102 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n16035), .ZN(P2_U3274) );
  AND2_X1 U17103 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n16035), .ZN(P2_U3273) );
  AND2_X1 U17104 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n16035), .ZN(P2_U3272) );
  AND2_X1 U17105 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n16035), .ZN(P2_U3271) );
  AND2_X1 U17106 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n16035), .ZN(P2_U3270) );
  AND2_X1 U17107 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n16035), .ZN(P2_U3269) );
  AND2_X1 U17108 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n16035), .ZN(P2_U3268) );
  AND2_X1 U17109 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n16035), .ZN(P2_U3267) );
  AND2_X1 U17110 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n16035), .ZN(P2_U3266) );
  NOR2_X1 U17111 ( .A1(n16110), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U17112 ( .A1(P3_U3897), .A2(n16036), .ZN(P3_U3150) );
  AOI22_X1 U17113 ( .A1(n16040), .A2(n16039), .B1(n16038), .B2(n16037), .ZN(
        P2_U3416) );
  AOI22_X1 U17114 ( .A1(n16110), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n16052) );
  OAI21_X1 U17115 ( .B1(n16043), .B2(n16042), .A(n16041), .ZN(n16044) );
  OAI22_X1 U17116 ( .A1(n16045), .A2(n16127), .B1(n16114), .B2(n16044), .ZN(
        n16046) );
  INV_X1 U17117 ( .A(n16046), .ZN(n16051) );
  OAI211_X1 U17118 ( .C1(n16049), .C2(n16048), .A(n16148), .B(n16047), .ZN(
        n16050) );
  NAND3_X1 U17119 ( .A1(n16052), .A2(n16051), .A3(n16050), .ZN(P2_U3215) );
  AOI22_X1 U17120 ( .A1(n16110), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n16064) );
  OAI21_X1 U17121 ( .B1(n16055), .B2(n16054), .A(n16053), .ZN(n16056) );
  OAI22_X1 U17122 ( .A1(n16057), .A2(n16127), .B1(n16114), .B2(n16056), .ZN(
        n16058) );
  INV_X1 U17123 ( .A(n16058), .ZN(n16063) );
  XOR2_X1 U17124 ( .A(n16060), .B(n16059), .Z(n16061) );
  NAND2_X1 U17125 ( .A1(n16148), .A2(n16061), .ZN(n16062) );
  NAND3_X1 U17126 ( .A1(n16064), .A2(n16063), .A3(n16062), .ZN(P2_U3216) );
  INV_X1 U17127 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n16203) );
  AND2_X1 U17128 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n16070) );
  OAI211_X1 U17129 ( .C1(n16067), .C2(n16066), .A(n16152), .B(n16065), .ZN(
        n16068) );
  INV_X1 U17130 ( .A(n16068), .ZN(n16069) );
  AOI211_X1 U17131 ( .C1(n16150), .C2(n16071), .A(n16070), .B(n16069), .ZN(
        n16076) );
  OAI211_X1 U17132 ( .C1(n16074), .C2(n16073), .A(n16148), .B(n16072), .ZN(
        n16075) );
  OAI211_X1 U17133 ( .C1(n16156), .C2(n16203), .A(n16076), .B(n16075), .ZN(
        P2_U3218) );
  AOI22_X1 U17134 ( .A1(n16110), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n16085) );
  OAI211_X1 U17135 ( .C1(n16078), .C2(P2_REG2_REG_15__SCAN_IN), .A(n16152), 
        .B(n16077), .ZN(n16084) );
  NAND2_X1 U17136 ( .A1(n16150), .A2(n16079), .ZN(n16083) );
  XNOR2_X1 U17137 ( .A(n16080), .B(P2_REG1_REG_15__SCAN_IN), .ZN(n16081) );
  NAND2_X1 U17138 ( .A1(n16081), .A2(n16148), .ZN(n16082) );
  NAND4_X1 U17139 ( .A1(n16085), .A2(n16084), .A3(n16083), .A4(n16082), .ZN(
        P2_U3229) );
  OAI21_X1 U17140 ( .B1(n16087), .B2(n16086), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n16088) );
  OAI21_X1 U17141 ( .B1(P2_STATE_REG_SCAN_IN), .B2(P2_REG3_REG_16__SCAN_IN), 
        .A(n16088), .ZN(n16098) );
  OAI211_X1 U17142 ( .C1(n16091), .C2(n16090), .A(n16089), .B(n16152), .ZN(
        n16097) );
  NAND2_X1 U17143 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n16110), .ZN(n16096) );
  OAI211_X1 U17144 ( .C1(n16094), .C2(n16093), .A(n16148), .B(n16092), .ZN(
        n16095) );
  NAND4_X1 U17145 ( .A1(n16098), .A2(n16097), .A3(n16096), .A4(n16095), .ZN(
        P2_U3230) );
  AOI22_X1 U17146 ( .A1(n16110), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3088), .ZN(n16109) );
  OAI211_X1 U17147 ( .C1(n16101), .C2(n16100), .A(n16152), .B(n16099), .ZN(
        n16108) );
  NAND2_X1 U17148 ( .A1(n16150), .A2(n16102), .ZN(n16107) );
  XOR2_X1 U17149 ( .A(n16104), .B(n16103), .Z(n16105) );
  NAND2_X1 U17150 ( .A1(n16148), .A2(n16105), .ZN(n16106) );
  NAND4_X1 U17151 ( .A1(n16109), .A2(n16108), .A3(n16107), .A4(n16106), .ZN(
        P2_U3231) );
  AOI22_X1 U17152 ( .A1(n16110), .A2(P2_ADDR_REG_18__SCAN_IN), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(P2_U3088), .ZN(n16121) );
  AOI21_X1 U17153 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n16112), .A(n16111), 
        .ZN(n16113) );
  OR2_X1 U17154 ( .A1(n16114), .A2(n16113), .ZN(n16120) );
  NAND2_X1 U17155 ( .A1(n16150), .A2(n16115), .ZN(n16119) );
  XOR2_X1 U17156 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n16116), .Z(n16117) );
  NAND2_X1 U17157 ( .A1(n16148), .A2(n16117), .ZN(n16118) );
  NAND4_X1 U17158 ( .A1(n16121), .A2(n16120), .A3(n16119), .A4(n16118), .ZN(
        P2_U3232) );
  INV_X1 U17159 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n16283) );
  NAND2_X1 U17160 ( .A1(n16123), .A2(n16122), .ZN(n16124) );
  NAND2_X1 U17161 ( .A1(n16125), .A2(n16124), .ZN(n16129) );
  NOR2_X1 U17162 ( .A1(n16127), .A2(n16126), .ZN(n16128) );
  AOI21_X1 U17163 ( .B1(n16129), .B2(n16148), .A(n16128), .ZN(n16136) );
  AND3_X1 U17164 ( .A1(n16132), .A2(n16131), .A3(n16130), .ZN(n16133) );
  OAI21_X1 U17165 ( .B1(n16134), .B2(n16133), .A(n16152), .ZN(n16135) );
  AND2_X1 U17166 ( .A1(n16136), .A2(n16135), .ZN(n16138) );
  OAI211_X1 U17167 ( .C1(n16283), .C2(n16156), .A(n16138), .B(n16137), .ZN(
        P2_U3226) );
  INV_X1 U17168 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n16157) );
  AND2_X1 U17169 ( .A1(n16140), .A2(n16139), .ZN(n16143) );
  OAI21_X1 U17170 ( .B1(n16143), .B2(n16142), .A(n16141), .ZN(n16153) );
  INV_X1 U17171 ( .A(n16144), .ZN(n16147) );
  MUX2_X1 U17172 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10302), .S(n16151), .Z(
        n16146) );
  OAI21_X1 U17173 ( .B1(n16147), .B2(n16146), .A(n16145), .ZN(n16149) );
  AOI222_X1 U17174 ( .A1(n16153), .A2(n16152), .B1(n16151), .B2(n16150), .C1(
        n16149), .C2(n16148), .ZN(n16155) );
  OAI211_X1 U17175 ( .C1(n16157), .C2(n16156), .A(n16155), .B(n16154), .ZN(
        P2_U3223) );
  OAI21_X1 U17176 ( .B1(n16159), .B2(P1_REG1_REG_0__SCAN_IN), .A(n16158), .ZN(
        n16161) );
  XNOR2_X1 U17177 ( .A(n16161), .B(n16160), .ZN(n16165) );
  AOI22_X1 U17178 ( .A1(n16162), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n16163) );
  OAI21_X1 U17179 ( .B1(n16165), .B2(n16164), .A(n16163), .ZN(P1_U3243) );
  INV_X1 U17180 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n16166) );
  AOI22_X1 U17181 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .B1(n16166), .B2(n16167), .ZN(n16168) );
  XOR2_X1 U17182 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n16168), .Z(SUB_1596_U53) );
  INV_X1 U17183 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n16180) );
  XOR2_X1 U17184 ( .A(n16172), .B(n16171), .Z(n16359) );
  NAND2_X1 U17185 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n16168), .ZN(n16358) );
  NAND2_X1 U17186 ( .A1(n16359), .A2(n16358), .ZN(n16169) );
  NOR2_X1 U17187 ( .A1(n16359), .A2(n16358), .ZN(n16357) );
  AOI21_X1 U17188 ( .B1(P2_ADDR_REG_1__SCAN_IN), .B2(n16169), .A(n16357), .ZN(
        n16170) );
  INV_X1 U17189 ( .A(n16170), .ZN(n16177) );
  NAND2_X1 U17190 ( .A1(n16172), .A2(n16171), .ZN(n16173) );
  XNOR2_X1 U17191 ( .A(n16175), .B(n16183), .ZN(n16185) );
  XNOR2_X1 U17192 ( .A(n16184), .B(n16185), .ZN(n16176) );
  NAND2_X1 U17193 ( .A1(n16177), .A2(n16176), .ZN(n16179) );
  NOR2_X1 U17194 ( .A1(n16177), .A2(n16176), .ZN(n16178) );
  INV_X1 U17195 ( .A(n16178), .ZN(n16182) );
  NAND2_X1 U17196 ( .A1(n16180), .A2(n16179), .ZN(n16181) );
  OAI222_X1 U17197 ( .A1(n16180), .A2(n16179), .B1(n16180), .B2(n16182), .C1(
        n16178), .C2(n16181), .ZN(SUB_1596_U61) );
  NAND2_X1 U17198 ( .A1(n16182), .A2(n16181), .ZN(n16197) );
  INV_X1 U17199 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n16188) );
  NAND2_X1 U17200 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n16183), .ZN(n16187) );
  NAND2_X1 U17201 ( .A1(n16185), .A2(n16184), .ZN(n16186) );
  NAND2_X1 U17202 ( .A1(n16187), .A2(n16186), .ZN(n16191) );
  XNOR2_X1 U17203 ( .A(n16188), .B(n16191), .ZN(n16193) );
  XNOR2_X1 U17204 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n16193), .ZN(n16198) );
  XOR2_X1 U17205 ( .A(n16197), .B(n16198), .Z(n16190) );
  INV_X1 U17206 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n16189) );
  NAND2_X1 U17207 ( .A1(n16190), .A2(n16189), .ZN(n16199) );
  OAI21_X1 U17208 ( .B1(n16190), .B2(n16189), .A(n16199), .ZN(SUB_1596_U60) );
  NAND2_X1 U17209 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n16191), .ZN(n16195) );
  NAND2_X1 U17210 ( .A1(n16193), .A2(n16192), .ZN(n16194) );
  NAND2_X1 U17211 ( .A1(n16195), .A2(n16194), .ZN(n16207) );
  XNOR2_X1 U17212 ( .A(n16196), .B(n16207), .ZN(n16209) );
  XNOR2_X1 U17213 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n16209), .ZN(n16204) );
  XNOR2_X1 U17214 ( .A(n16203), .B(n16204), .ZN(n16202) );
  NAND2_X1 U17215 ( .A1(n16198), .A2(n16197), .ZN(n16200) );
  NAND2_X1 U17216 ( .A1(n16200), .A2(n16199), .ZN(n16201) );
  NOR2_X1 U17217 ( .A1(n16202), .A2(n16201), .ZN(n16205) );
  AOI21_X1 U17218 ( .B1(n16202), .B2(n16201), .A(n16205), .ZN(SUB_1596_U59) );
  NOR2_X1 U17219 ( .A1(n16204), .A2(n16203), .ZN(n16206) );
  NAND2_X1 U17220 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n16207), .ZN(n16211) );
  NAND2_X1 U17221 ( .A1(n16209), .A2(n16208), .ZN(n16210) );
  NAND2_X1 U17222 ( .A1(n16211), .A2(n16210), .ZN(n16214) );
  NOR2_X1 U17223 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n16217), .ZN(n16212) );
  AOI21_X1 U17224 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(n16217), .A(n16212), .ZN(
        n16215) );
  XOR2_X1 U17225 ( .A(n16214), .B(n16215), .Z(n16219) );
  NAND2_X1 U17226 ( .A1(n16220), .A2(n16219), .ZN(n16221) );
  OAI21_X1 U17227 ( .B1(n16220), .B2(n16219), .A(n16221), .ZN(n16213) );
  XNOR2_X1 U17228 ( .A(n16213), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  NAND2_X1 U17229 ( .A1(n16215), .A2(n16214), .ZN(n16216) );
  XOR2_X1 U17230 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), .Z(
        n16218) );
  XNOR2_X1 U17231 ( .A(n16225), .B(n16218), .ZN(n16355) );
  NAND2_X1 U17232 ( .A1(n16355), .A2(n16354), .ZN(n16353) );
  XNOR2_X1 U17233 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n16235), .ZN(n16228) );
  INV_X1 U17234 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n16230) );
  INV_X1 U17235 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n16223) );
  NOR2_X1 U17236 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n16223), .ZN(n16226) );
  NAND2_X1 U17237 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n16223), .ZN(n16224) );
  XNOR2_X1 U17238 ( .A(n16230), .B(n16229), .ZN(n16231) );
  XOR2_X1 U17239 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n16231), .Z(n16227) );
  NAND2_X1 U17240 ( .A1(n16228), .A2(n16227), .ZN(n16237) );
  OAI21_X1 U17241 ( .B1(n16228), .B2(n16227), .A(n16237), .ZN(SUB_1596_U56) );
  INV_X1 U17242 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n16243) );
  NOR2_X1 U17243 ( .A1(n16230), .A2(n16229), .ZN(n16233) );
  AOI22_X1 U17244 ( .A1(P3_ADDR_REG_8__SCAN_IN), .A2(n16234), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n16246), .ZN(n16248) );
  XOR2_X1 U17245 ( .A(n16247), .B(n16248), .Z(n16240) );
  INV_X1 U17246 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n16236) );
  NAND2_X1 U17247 ( .A1(n16236), .A2(n16235), .ZN(n16238) );
  AND2_X2 U17248 ( .A1(n16238), .A2(n16237), .ZN(n16239) );
  NAND2_X1 U17249 ( .A1(n16240), .A2(n16239), .ZN(n16242) );
  NAND2_X1 U17250 ( .A1(n16243), .A2(n16242), .ZN(n16244) );
  OAI222_X1 U17251 ( .A1(n16243), .A2(n16242), .B1(n16243), .B2(n16245), .C1(
        n16241), .C2(n16244), .ZN(SUB_1596_U55) );
  NAND2_X1 U17252 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n16246), .ZN(n16250) );
  NAND2_X1 U17253 ( .A1(n16248), .A2(n16247), .ZN(n16249) );
  NAND2_X1 U17254 ( .A1(n16250), .A2(n16249), .ZN(n16258) );
  AOI22_X1 U17255 ( .A1(P3_ADDR_REG_9__SCAN_IN), .A2(n16251), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n16257), .ZN(n16259) );
  XNOR2_X1 U17256 ( .A(n16258), .B(n16259), .ZN(n16253) );
  AOI21_X1 U17257 ( .B1(n16254), .B2(n16253), .A(n16255), .ZN(n16252) );
  XOR2_X1 U17258 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n16252), .Z(SUB_1596_U54) );
  NAND2_X1 U17259 ( .A1(n16254), .A2(n16253), .ZN(n16256) );
  NAND2_X1 U17260 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n16257), .ZN(n16261) );
  NAND2_X1 U17261 ( .A1(n16259), .A2(n16258), .ZN(n16260) );
  NAND2_X1 U17262 ( .A1(n16261), .A2(n16260), .ZN(n16264) );
  XOR2_X1 U17263 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n16263) );
  XOR2_X1 U17264 ( .A(n16264), .B(n16263), .Z(n16267) );
  NAND2_X1 U17265 ( .A1(n16268), .A2(n16267), .ZN(n16269) );
  OAI21_X1 U17266 ( .B1(n16268), .B2(n16267), .A(n16269), .ZN(n16262) );
  XNOR2_X1 U17267 ( .A(n16262), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  INV_X1 U17268 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n16276) );
  INV_X1 U17269 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n16282) );
  XNOR2_X1 U17270 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(n16282), .ZN(n16280) );
  INV_X1 U17271 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n16266) );
  XOR2_X1 U17272 ( .A(n16280), .B(n16279), .Z(n16273) );
  NOR2_X1 U17273 ( .A1(n16268), .A2(n16267), .ZN(n16270) );
  OAI21_X1 U17274 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(n16270), .A(n16269), 
        .ZN(n16271) );
  INV_X1 U17275 ( .A(n16271), .ZN(n16272) );
  NAND2_X1 U17276 ( .A1(n16273), .A2(n16272), .ZN(n16275) );
  NAND2_X1 U17277 ( .A1(n16276), .A2(n16275), .ZN(n16277) );
  OAI222_X1 U17278 ( .A1(n16276), .A2(n16275), .B1(n16276), .B2(n16278), .C1(
        n16274), .C2(n16277), .ZN(SUB_1596_U69) );
  XOR2_X1 U17279 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .Z(n16285) );
  XOR2_X1 U17280 ( .A(n16286), .B(n16285), .Z(n16291) );
  NAND2_X1 U17281 ( .A1(n16284), .A2(n16283), .ZN(n16292) );
  OAI21_X1 U17282 ( .B1(n16284), .B2(n16283), .A(n16292), .ZN(SUB_1596_U68) );
  XOR2_X1 U17283 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n16289) );
  XOR2_X1 U17284 ( .A(n16301), .B(n16289), .Z(n16296) );
  NAND2_X1 U17285 ( .A1(n16291), .A2(n16290), .ZN(n16293) );
  NAND2_X1 U17286 ( .A1(n16296), .A2(n16295), .ZN(n16297) );
  OAI21_X1 U17287 ( .B1(n16296), .B2(n16295), .A(n16297), .ZN(n16294) );
  XNOR2_X1 U17288 ( .A(n16294), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  NOR2_X1 U17289 ( .A1(n16296), .A2(n16295), .ZN(n16298) );
  INV_X1 U17290 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n16302) );
  INV_X1 U17291 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n16299) );
  NOR2_X1 U17292 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n16299), .ZN(n16300) );
  XNOR2_X1 U17293 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n16308) );
  XOR2_X1 U17294 ( .A(n16307), .B(n16308), .Z(n16305) );
  OAI21_X1 U17295 ( .B1(n16304), .B2(n16305), .A(n16306), .ZN(n16303) );
  XNOR2_X1 U17296 ( .A(n16303), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  XNOR2_X1 U17297 ( .A(P3_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n16311) );
  INV_X1 U17298 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n16310) );
  NAND2_X1 U17299 ( .A1(n16308), .A2(n16307), .ZN(n16309) );
  XOR2_X1 U17300 ( .A(n16311), .B(n16314), .Z(n16316) );
  AOI21_X1 U17301 ( .B1(n16317), .B2(n16316), .A(n16318), .ZN(n16312) );
  XOR2_X1 U17302 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n16312), .Z(SUB_1596_U65)
         );
  INV_X1 U17303 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n16365) );
  NAND2_X1 U17304 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n16365), .ZN(n16313) );
  AOI22_X1 U17305 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n16315), .B1(n16314), 
        .B2(n16313), .ZN(n16325) );
  XOR2_X1 U17306 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n16325), .Z(n16327) );
  XNOR2_X1 U17307 ( .A(n16326), .B(n16327), .ZN(n16321) );
  NAND2_X1 U17308 ( .A1(n16317), .A2(n16316), .ZN(n16319) );
  NAND2_X1 U17309 ( .A1(n16322), .A2(n16321), .ZN(n16323) );
  OAI21_X1 U17310 ( .B1(n16321), .B2(n16322), .A(n16323), .ZN(n16320) );
  XNOR2_X1 U17311 ( .A(n16320), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  NOR2_X1 U17312 ( .A1(n16322), .A2(n16321), .ZN(n16324) );
  OAI21_X1 U17313 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(n16324), .A(n16323), 
        .ZN(n16331) );
  NAND2_X1 U17314 ( .A1(n16325), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n16329) );
  NAND2_X1 U17315 ( .A1(n16327), .A2(n16326), .ZN(n16328) );
  NAND2_X1 U17316 ( .A1(n16329), .A2(n16328), .ZN(n16335) );
  XNOR2_X1 U17317 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n16335), .ZN(n16336) );
  XOR2_X1 U17318 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n16336), .Z(n16332) );
  XNOR2_X1 U17319 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n16332), .ZN(n16330) );
  NOR2_X1 U17320 ( .A1(n16331), .A2(n16330), .ZN(n16333) );
  AOI21_X1 U17321 ( .B1(n16331), .B2(n16330), .A(n16333), .ZN(SUB_1596_U63) );
  AND2_X1 U17322 ( .A1(n16332), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n16334) );
  NOR2_X1 U17323 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n16335), .ZN(n16339) );
  INV_X1 U17324 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n16337) );
  NOR2_X1 U17325 ( .A1(n16337), .A2(n16336), .ZN(n16338) );
  NOR2_X1 U17326 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n16345), .ZN(n16340) );
  AOI21_X1 U17327 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n16345), .A(n16340), 
        .ZN(n16343) );
  XOR2_X1 U17328 ( .A(n16342), .B(n16343), .Z(n16346) );
  OAI21_X1 U17329 ( .B1(n16347), .B2(n16346), .A(n16348), .ZN(n16341) );
  XNOR2_X1 U17330 ( .A(n16341), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NAND2_X1 U17331 ( .A1(n16343), .A2(n16342), .ZN(n16344) );
  OAI21_X1 U17332 ( .B1(n16345), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n16344), 
        .ZN(n16352) );
  XNOR2_X1 U17333 ( .A(n16349), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n16350) );
  XNOR2_X1 U17334 ( .A(n16350), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n16351) );
  OAI21_X1 U17335 ( .B1(n16355), .B2(n16354), .A(n16353), .ZN(n16356) );
  XNOR2_X1 U17336 ( .A(n16356), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(SUB_1596_U57)
         );
  AOI21_X1 U17337 ( .B1(n16359), .B2(n16358), .A(n16357), .ZN(n16360) );
  XOR2_X1 U17338 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n16360), .Z(SUB_1596_U5) );
  AOI21_X1 U17339 ( .B1(n16363), .B2(n16362), .A(n16361), .ZN(n16383) );
  OAI22_X1 U17340 ( .A1(n16367), .A2(n16366), .B1(n16365), .B2(n16364), .ZN(
        n16379) );
  AOI21_X1 U17341 ( .B1(n16370), .B2(n16369), .A(n16368), .ZN(n16377) );
  AOI21_X1 U17342 ( .B1(n16373), .B2(n16372), .A(n16371), .ZN(n16375) );
  OAI22_X1 U17343 ( .A1(n16377), .A2(n16376), .B1(n16375), .B2(n16374), .ZN(
        n16378) );
  NOR3_X1 U17344 ( .A1(n16380), .A2(n16379), .A3(n16378), .ZN(n16381) );
  OAI21_X1 U17345 ( .B1(n16383), .B2(n16382), .A(n16381), .ZN(P3_U3197) );
  OAI221_X1 U17346 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(
        n16385), .C2(n8434), .A(n16384), .ZN(U29) );
  INV_X1 U17347 ( .A(n16493), .ZN(n16412) );
  AND2_X1 U17348 ( .A1(n16386), .A2(n8315), .ZN(n16393) );
  OAI21_X1 U17349 ( .B1(n16387), .B2(n16458), .A(n16398), .ZN(n16388) );
  OAI21_X1 U17350 ( .B1(n7600), .B2(n16389), .A(n16388), .ZN(n16396) );
  AOI211_X1 U17351 ( .C1(n16412), .C2(n16398), .A(n16393), .B(n16396), .ZN(
        n16391) );
  AOI22_X1 U17352 ( .A1(n16469), .A2(n16391), .B1(n16390), .B2(n16565), .ZN(
        P1_U3528) );
  AOI22_X1 U17353 ( .A1(n16570), .A2(n16391), .B1(n10351), .B2(n16567), .ZN(
        P1_U3459) );
  NAND2_X1 U17354 ( .A1(n16393), .A2(n16392), .ZN(n16394) );
  OAI21_X1 U17355 ( .B1(n16395), .B2(n10349), .A(n16394), .ZN(n16397) );
  AOI211_X1 U17356 ( .C1(n16399), .C2(n16398), .A(n16397), .B(n16396), .ZN(
        n16400) );
  AOI22_X1 U17357 ( .A1(n16605), .A2(n16401), .B1(n16400), .B2(n15812), .ZN(
        P1_U3293) );
  AOI211_X1 U17358 ( .C1(n16578), .C2(n16404), .A(n16403), .B(n16402), .ZN(
        n16406) );
  AOI22_X1 U17359 ( .A1(n16587), .A2(n16406), .B1(n16405), .B2(n16585), .ZN(
        P3_U3460) );
  AOI22_X1 U17360 ( .A1(n16590), .A2(n16406), .B1(n9599), .B2(n16588), .ZN(
        P3_U3393) );
  OAI21_X1 U17361 ( .B1(n7601), .B2(n16556), .A(n16407), .ZN(n16410) );
  INV_X1 U17362 ( .A(n16408), .ZN(n16409) );
  AOI211_X1 U17363 ( .C1(n16412), .C2(n16411), .A(n16410), .B(n16409), .ZN(
        n16415) );
  AOI22_X1 U17364 ( .A1(n16469), .A2(n16415), .B1(n16413), .B2(n16565), .ZN(
        P1_U3529) );
  INV_X1 U17365 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n16414) );
  AOI22_X1 U17366 ( .A1(n16570), .A2(n16415), .B1(n16414), .B2(n16567), .ZN(
        P1_U3462) );
  AOI22_X1 U17367 ( .A1(P2_REG2_REG_1__SCAN_IN), .A2(n16522), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n16511), .ZN(n16422) );
  AOI222_X1 U17368 ( .A1(n16420), .A2(n16419), .B1(n16418), .B2(n16508), .C1(
        n16417), .C2(n16416), .ZN(n16421) );
  OAI211_X1 U17369 ( .C1(n16522), .C2(n16423), .A(n16422), .B(n16421), .ZN(
        P2_U3264) );
  INV_X1 U17370 ( .A(n16424), .ZN(n16426) );
  AOI211_X1 U17371 ( .C1(n16485), .C2(n16427), .A(n16426), .B(n16425), .ZN(
        n16430) );
  AOI22_X1 U17372 ( .A1(n16587), .A2(n16430), .B1(n16428), .B2(n16585), .ZN(
        P3_U3461) );
  INV_X1 U17373 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n16429) );
  AOI22_X1 U17374 ( .A1(n16590), .A2(n16430), .B1(n16429), .B2(n16588), .ZN(
        P3_U3396) );
  INV_X1 U17375 ( .A(n16431), .ZN(n16433) );
  OAI211_X1 U17376 ( .C1(n16434), .C2(n16556), .A(n16433), .B(n16432), .ZN(
        n16438) );
  NOR2_X1 U17377 ( .A1(n16436), .A2(n16435), .ZN(n16437) );
  AOI211_X1 U17378 ( .C1(n16458), .C2(n16439), .A(n16438), .B(n16437), .ZN(
        n16442) );
  AOI22_X1 U17379 ( .A1(n16469), .A2(n16442), .B1(n16440), .B2(n16565), .ZN(
        P1_U3530) );
  INV_X1 U17380 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n16441) );
  AOI22_X1 U17381 ( .A1(n16570), .A2(n16442), .B1(n16441), .B2(n16567), .ZN(
        P1_U3465) );
  AOI22_X1 U17382 ( .A1(n15102), .A2(n16443), .B1(n8573), .B2(n16623), .ZN(
        P2_U3436) );
  NOR2_X1 U17383 ( .A1(n16444), .A2(n16580), .ZN(n16446) );
  AOI211_X1 U17384 ( .C1(n16485), .C2(n16447), .A(n16446), .B(n16445), .ZN(
        n16449) );
  AOI22_X1 U17385 ( .A1(n16587), .A2(n16449), .B1(n16448), .B2(n16585), .ZN(
        P3_U3462) );
  AOI22_X1 U17386 ( .A1(n16590), .A2(n16449), .B1(n9620), .B2(n16588), .ZN(
        P3_U3399) );
  OAI211_X1 U17387 ( .C1(n16452), .C2(n16556), .A(n16451), .B(n16450), .ZN(
        n16456) );
  AOI21_X1 U17388 ( .B1(n16493), .B2(n16454), .A(n16453), .ZN(n16455) );
  AOI211_X1 U17389 ( .C1(n16458), .C2(n16457), .A(n16456), .B(n16455), .ZN(
        n16460) );
  AOI22_X1 U17390 ( .A1(n16469), .A2(n16460), .B1(n10504), .B2(n16565), .ZN(
        P1_U3531) );
  INV_X1 U17391 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n16459) );
  AOI22_X1 U17392 ( .A1(n16570), .A2(n16460), .B1(n16459), .B2(n16567), .ZN(
        P1_U3468) );
  INV_X1 U17393 ( .A(n16461), .ZN(n16462) );
  OAI21_X1 U17394 ( .B1(n16463), .B2(n16556), .A(n16462), .ZN(n16466) );
  INV_X1 U17395 ( .A(n16464), .ZN(n16465) );
  AOI211_X1 U17396 ( .C1(n16467), .C2(n16564), .A(n16466), .B(n16465), .ZN(
        n16471) );
  AOI22_X1 U17397 ( .A1(n16469), .A2(n16471), .B1(n16468), .B2(n16565), .ZN(
        P1_U3532) );
  INV_X1 U17398 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n16470) );
  AOI22_X1 U17399 ( .A1(n16570), .A2(n16471), .B1(n16470), .B2(n16567), .ZN(
        P1_U3471) );
  INV_X1 U17400 ( .A(n16472), .ZN(n16473) );
  AOI22_X1 U17401 ( .A1(n14992), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n16473), 
        .B2(n16511), .ZN(n16474) );
  OAI21_X1 U17402 ( .B1(n16515), .B2(n16475), .A(n16474), .ZN(n16476) );
  INV_X1 U17403 ( .A(n16476), .ZN(n16480) );
  AOI22_X1 U17404 ( .A1(n16519), .A2(n16478), .B1(n16508), .B2(n16477), .ZN(
        n16479) );
  OAI211_X1 U17405 ( .C1(n16522), .C2(n16481), .A(n16480), .B(n16479), .ZN(
        P2_U3261) );
  NOR2_X1 U17406 ( .A1(n9997), .A2(n16580), .ZN(n16483) );
  AOI211_X1 U17407 ( .C1(n16485), .C2(n16484), .A(n16483), .B(n16482), .ZN(
        n16487) );
  AOI22_X1 U17408 ( .A1(n16587), .A2(n16487), .B1(n16486), .B2(n16585), .ZN(
        P3_U3464) );
  AOI22_X1 U17409 ( .A1(n16590), .A2(n16487), .B1(n9650), .B2(n16588), .ZN(
        P3_U3405) );
  AOI21_X1 U17410 ( .B1(n16490), .B2(n16489), .A(n16488), .ZN(n16491) );
  OAI211_X1 U17411 ( .C1(n16494), .C2(n16493), .A(n16492), .B(n16491), .ZN(
        n16495) );
  INV_X1 U17412 ( .A(n16495), .ZN(n16497) );
  AOI22_X1 U17413 ( .A1(n16469), .A2(n16497), .B1(n16496), .B2(n16565), .ZN(
        P1_U3534) );
  AOI22_X1 U17414 ( .A1(n16570), .A2(n16497), .B1(n10801), .B2(n16567), .ZN(
        P1_U3477) );
  OAI21_X1 U17415 ( .B1(n16499), .B2(n16616), .A(n16498), .ZN(n16501) );
  AOI211_X1 U17416 ( .C1(n16610), .C2(n16502), .A(n16501), .B(n16500), .ZN(
        n16504) );
  AOI22_X1 U17417 ( .A1(n7433), .A2(n16504), .B1(n10292), .B2(n16622), .ZN(
        P2_U3505) );
  INV_X1 U17418 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n16503) );
  AOI22_X1 U17419 ( .A1(n15102), .A2(n16504), .B1(n16503), .B2(n16623), .ZN(
        P2_U3448) );
  INV_X1 U17420 ( .A(n16505), .ZN(n16506) );
  AOI21_X1 U17421 ( .B1(n16507), .B2(n16518), .A(n16506), .ZN(n16521) );
  NAND2_X1 U17422 ( .A1(n16509), .A2(n16508), .ZN(n16514) );
  INV_X1 U17423 ( .A(n16510), .ZN(n16512) );
  AOI22_X1 U17424 ( .A1(n14992), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n16512), 
        .B2(n16511), .ZN(n16513) );
  OAI211_X1 U17425 ( .C1(n16516), .C2(n16515), .A(n16514), .B(n16513), .ZN(
        n16517) );
  AOI21_X1 U17426 ( .B1(n16519), .B2(n16518), .A(n16517), .ZN(n16520) );
  OAI21_X1 U17427 ( .B1(n16522), .B2(n16521), .A(n16520), .ZN(P2_U3258) );
  INV_X1 U17428 ( .A(n16523), .ZN(n16524) );
  AOI222_X1 U17429 ( .A1(n16526), .A2(n16525), .B1(n16524), .B2(n16592), .C1(
        P1_REG2_REG_8__SCAN_IN), .C2(n16605), .ZN(n16531) );
  INV_X1 U17430 ( .A(n16547), .ZN(n16528) );
  AOI22_X1 U17431 ( .A1(n16529), .A2(n16528), .B1(n16601), .B2(n16527), .ZN(
        n16530) );
  OAI211_X1 U17432 ( .C1(n16605), .C2(n16532), .A(n16531), .B(n16530), .ZN(
        P1_U3285) );
  OAI21_X1 U17433 ( .B1(n7947), .B2(n16616), .A(n16533), .ZN(n16535) );
  AOI211_X1 U17434 ( .C1(n16536), .C2(n16621), .A(n16535), .B(n16534), .ZN(
        n16537) );
  AOI22_X1 U17435 ( .A1(n7433), .A2(n16537), .B1(n10298), .B2(n16622), .ZN(
        P2_U3507) );
  AOI22_X1 U17436 ( .A1(n15102), .A2(n16537), .B1(n8721), .B2(n16623), .ZN(
        P2_U3454) );
  AOI22_X1 U17437 ( .A1(n16540), .A2(n16587), .B1(n16539), .B2(n16538), .ZN(
        n16541) );
  OAI21_X1 U17438 ( .B1(n16587), .B2(n16542), .A(n16541), .ZN(P3_U3468) );
  INV_X1 U17439 ( .A(n16543), .ZN(n16544) );
  AOI22_X1 U17440 ( .A1(n16605), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n16544), 
        .B2(n16592), .ZN(n16545) );
  OAI21_X1 U17441 ( .B1(n16546), .B2(n16595), .A(n16545), .ZN(n16550) );
  NOR2_X1 U17442 ( .A1(n16548), .A2(n16547), .ZN(n16549) );
  AOI211_X1 U17443 ( .C1(n16551), .C2(n16601), .A(n16550), .B(n16549), .ZN(
        n16552) );
  OAI21_X1 U17444 ( .B1(n16605), .B2(n16553), .A(n16552), .ZN(P1_U3284) );
  OAI211_X1 U17445 ( .C1(n16557), .C2(n16556), .A(n16555), .B(n16554), .ZN(
        n16562) );
  NOR3_X1 U17446 ( .A1(n16560), .A2(n16559), .A3(n16558), .ZN(n16561) );
  AOI211_X1 U17447 ( .C1(n16564), .C2(n16563), .A(n16562), .B(n16561), .ZN(
        n16569) );
  AOI22_X1 U17448 ( .A1(n16469), .A2(n16569), .B1(n16566), .B2(n16565), .ZN(
        P1_U3538) );
  INV_X1 U17449 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n16568) );
  AOI22_X1 U17450 ( .A1(n16570), .A2(n16569), .B1(n16568), .B2(n16567), .ZN(
        P1_U3489) );
  OAI211_X1 U17451 ( .C1(n16573), .C2(n16616), .A(n16572), .B(n16571), .ZN(
        n16574) );
  AOI21_X1 U17452 ( .B1(n16621), .B2(n16575), .A(n16574), .ZN(n16577) );
  AOI22_X1 U17453 ( .A1(n7433), .A2(n16577), .B1(n16576), .B2(n16622), .ZN(
        P2_U3509) );
  AOI22_X1 U17454 ( .A1(n15102), .A2(n16577), .B1(n8758), .B2(n16623), .ZN(
        P2_U3460) );
  AND2_X1 U17455 ( .A1(n16579), .A2(n16578), .ZN(n16584) );
  NOR2_X1 U17456 ( .A1(n16581), .A2(n16580), .ZN(n16583) );
  NOR3_X1 U17457 ( .A1(n16584), .A2(n16583), .A3(n16582), .ZN(n16589) );
  AOI22_X1 U17458 ( .A1(n16587), .A2(n16589), .B1(n16586), .B2(n16585), .ZN(
        P3_U3470) );
  AOI22_X1 U17459 ( .A1(n16590), .A2(n16589), .B1(n9738), .B2(n16588), .ZN(
        P3_U3423) );
  INV_X1 U17460 ( .A(n16591), .ZN(n16593) );
  AOI22_X1 U17461 ( .A1(n16605), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n16593), 
        .B2(n16592), .ZN(n16594) );
  OAI21_X1 U17462 ( .B1(n16596), .B2(n16595), .A(n16594), .ZN(n16600) );
  NOR2_X1 U17463 ( .A1(n16598), .A2(n16597), .ZN(n16599) );
  AOI211_X1 U17464 ( .C1(n16602), .C2(n16601), .A(n16600), .B(n16599), .ZN(
        n16603) );
  OAI21_X1 U17465 ( .B1(n16605), .B2(n16604), .A(n16603), .ZN(P1_U3282) );
  INV_X1 U17466 ( .A(n16606), .ZN(n16608) );
  OAI21_X1 U17467 ( .B1(n16608), .B2(n16616), .A(n16607), .ZN(n16609) );
  AOI21_X1 U17468 ( .B1(n16611), .B2(n16610), .A(n16609), .ZN(n16612) );
  AND2_X1 U17469 ( .A1(n16613), .A2(n16612), .ZN(n16614) );
  AOI22_X1 U17470 ( .A1(n7433), .A2(n16614), .B1(n10569), .B2(n16622), .ZN(
        P2_U3511) );
  AOI22_X1 U17471 ( .A1(n15102), .A2(n16614), .B1(n8806), .B2(n16623), .ZN(
        P2_U3466) );
  OAI21_X1 U17472 ( .B1(n16617), .B2(n16616), .A(n16615), .ZN(n16619) );
  AOI211_X1 U17473 ( .C1(n16621), .C2(n16620), .A(n16619), .B(n16618), .ZN(
        n16624) );
  AOI22_X1 U17474 ( .A1(n7433), .A2(n16624), .B1(n8839), .B2(n16622), .ZN(
        P2_U3513) );
  AOI22_X1 U17475 ( .A1(n15102), .A2(n16624), .B1(n8840), .B2(n16623), .ZN(
        P2_U3472) );
  AOI21_X1 U17476 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16625) );
  OAI21_X1 U17477 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16625), 
        .ZN(U28) );
  AND3_X1 U7583 ( .A1(n9588), .A2(n9587), .A3(n9589), .ZN(n9591) );
  CLKBUF_X1 U7542 ( .A(n7604), .Z(n7427) );
  CLKBUF_X1 U7555 ( .A(n8969), .Z(n9341) );
  AOI21_X2 U7597 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(n16319), .A(n16318), .ZN(
        n16322) );
endmodule

