

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n5081, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11044;

  CLKBUF_X2 U5145 ( .A(n6681), .Z(n6956) );
  INV_X1 U5146 ( .A(n5084), .ZN(n5085) );
  AND2_X1 U5147 ( .A1(n10584), .A2(n8790), .ZN(n6667) );
  NAND2_X1 U5148 ( .A1(n5597), .A2(n5595), .ZN(n5974) );
  NOR2_X1 U5149 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5504) );
  INV_X1 U5150 ( .A(n11044), .ZN(n5081) );
  INV_X2 U5151 ( .A(n5081), .ZN(P2_U3151) );
  INV_X1 U5152 ( .A(P2_STATE_REG_SCAN_IN), .ZN(n11044) );
  NAND2_X2 U5153 ( .A1(n10574), .A2(n10573), .ZN(n10590) );
  OAI21_X1 U5154 ( .B1(n7441), .B2(n5819), .A(n7491), .ZN(n5307) );
  NAND2_X1 U5155 ( .A1(n5780), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5777) );
  INV_X2 U5156 ( .A(n9951), .ZN(n9899) );
  INV_X1 U5157 ( .A(n7735), .ZN(n7766) );
  INV_X1 U5158 ( .A(n6128), .ZN(n7312) );
  OAI21_X1 U5159 ( .B1(n9496), .B2(n5499), .A(n5498), .ZN(n5895) );
  CLKBUF_X3 U5160 ( .A(n6085), .Z(n7301) );
  AND2_X1 U5161 ( .A1(n5450), .A2(n7511), .ZN(n9953) );
  INV_X1 U5162 ( .A(n8072), .ZN(n10838) );
  INV_X2 U5163 ( .A(n7808), .ZN(n9863) );
  INV_X2 U5164 ( .A(n6682), .ZN(n6794) );
  NAND2_X1 U5165 ( .A1(n7151), .A2(n7150), .ZN(n7410) );
  INV_X1 U5166 ( .A(n8034), .ZN(n7806) );
  AND4_X1 U5167 ( .A1(n5964), .A2(n5963), .A3(n5962), .A4(n5961), .ZN(n9589)
         );
  AND4_X1 U5168 ( .A1(n6426), .A2(n6425), .A3(n6424), .A4(n6423), .ZN(n10659)
         );
  AND3_X1 U5169 ( .A1(n5803), .A2(n5735), .A3(n5736), .ZN(n5083) );
  NOR2_X2 U5170 ( .A1(n7152), .A2(n6559), .ZN(n6560) );
  OR2_X2 U5171 ( .A1(n9403), .A2(n7930), .ZN(n7191) );
  NAND2_X2 U5172 ( .A1(n6679), .A2(n7081), .ZN(n10783) );
  AOI21_X2 U5173 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n7374), .A(n7454), .ZN(
        n5877) );
  AND2_X1 U5174 ( .A1(n6574), .A2(n8790), .ZN(n5091) );
  AOI21_X2 U5175 ( .B1(n10316), .B2(n10244), .A(n10243), .ZN(n10303) );
  NAND2_X2 U5176 ( .A1(n10333), .A2(n10242), .ZN(n10316) );
  INV_X1 U5177 ( .A(n7363), .ZN(n7450) );
  NOR2_X2 U5178 ( .A1(n6167), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6182) );
  XNOR2_X2 U5179 ( .A(n6556), .B(n9236), .ZN(n7150) );
  NAND2_X4 U5180 ( .A1(n9259), .A2(n9256), .ZN(n6470) );
  XNOR2_X2 U5181 ( .A(n5777), .B(n5951), .ZN(n5864) );
  NOR2_X2 U5182 ( .A1(n7443), .A2(n7442), .ZN(n7441) );
  INV_X2 U5183 ( .A(n6116), .ZN(n5084) );
  INV_X4 U5184 ( .A(n5084), .ZN(n5086) );
  NAND2_X1 U5185 ( .A1(n9259), .A2(n5958), .ZN(n6116) );
  XNOR2_X2 U5186 ( .A(n5884), .B(n8505), .ZN(n8496) );
  NOR2_X2 U5187 ( .A1(n8198), .A2(n5883), .ZN(n5884) );
  AND2_X1 U5188 ( .A1(n6386), .A2(n9296), .ZN(n6388) );
  NAND2_X1 U5189 ( .A1(n10101), .A2(n10838), .ZN(n7086) );
  NAND2_X1 U5190 ( .A1(n7084), .A2(n7000), .ZN(n8032) );
  NAND2_X1 U5191 ( .A1(n8011), .A2(n7046), .ZN(n10818) );
  INV_X1 U5192 ( .A(n10829), .ZN(n10816) );
  INV_X1 U5193 ( .A(n7772), .ZN(n8312) );
  INV_X2 U5194 ( .A(n7754), .ZN(n8401) );
  INV_X1 U5195 ( .A(n7547), .ZN(n6976) );
  OAI21_X1 U5196 ( .B1(n9912), .B2(n9959), .A(n10081), .ZN(n9917) );
  OAI21_X1 U5197 ( .B1(n9983), .B2(n5282), .A(n5279), .ZN(n9958) );
  NAND2_X1 U5198 ( .A1(n9918), .A2(n5443), .ZN(n5445) );
  AND2_X1 U5199 ( .A1(n9814), .A2(n5178), .ZN(n5443) );
  NAND2_X1 U5200 ( .A1(n9263), .A2(n9622), .ZN(n9262) );
  OR2_X1 U5201 ( .A1(n5296), .A2(n5153), .ZN(n5294) );
  XNOR2_X1 U5202 ( .A(n8824), .B(n8825), .ZN(n9263) );
  NOR2_X1 U5203 ( .A1(n9811), .A2(n9810), .ZN(n9813) );
  NOR2_X1 U5204 ( .A1(n9497), .A2(n9498), .ZN(n9496) );
  OR2_X1 U5205 ( .A1(n5892), .A2(n5894), .ZN(n5499) );
  XNOR2_X1 U5206 ( .A(n9584), .B(n9386), .ZN(n9579) );
  NAND2_X1 U5207 ( .A1(n5350), .A2(n5348), .ZN(n6460) );
  NOR2_X1 U5208 ( .A1(n9488), .A2(n5714), .ZN(n5859) );
  XNOR2_X1 U5209 ( .A(n6393), .B(n9387), .ZN(n9594) );
  OAI21_X1 U5210 ( .B1(n8299), .B2(n8298), .A(n8297), .ZN(n8301) );
  NAND2_X1 U5211 ( .A1(n8558), .A2(n8557), .ZN(n8636) );
  AOI21_X1 U5212 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n9449), .A(n9450), .ZN(
        n5849) );
  NAND2_X1 U5213 ( .A1(n8068), .A2(n8067), .ZN(n8147) );
  NAND2_X1 U5214 ( .A1(n8065), .A2(n8064), .ZN(n8070) );
  NAND2_X1 U5215 ( .A1(n5447), .A2(n5244), .ZN(n8065) );
  OAI21_X1 U5216 ( .B1(n6358), .B2(n6357), .A(n6046), .ZN(n6064) );
  OAI21_X1 U5217 ( .B1(n7009), .B2(n5526), .A(n5524), .ZN(n10946) );
  NAND2_X1 U5218 ( .A1(n7825), .A2(n7824), .ZN(n5447) );
  OR2_X1 U5219 ( .A1(n9416), .A2(n5886), .ZN(n5888) );
  OAI21_X1 U5220 ( .B1(n6026), .B2(n5590), .A(n5588), .ZN(n6333) );
  NAND2_X1 U5221 ( .A1(n6852), .A2(n6851), .ZN(n10556) );
  NOR2_X1 U5222 ( .A1(n5448), .A2(n7839), .ZN(n5244) );
  NAND2_X1 U5223 ( .A1(n6811), .A2(n6810), .ZN(n10957) );
  INV_X1 U5224 ( .A(n6419), .ZN(n6406) );
  NOR2_X1 U5225 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(n6419), .ZN(n6420) );
  NAND2_X1 U5226 ( .A1(n6388), .A2(n9375), .ZN(n6419) );
  NAND2_X1 U5227 ( .A1(n6790), .A2(n6789), .ZN(n8619) );
  AND2_X1 U5228 ( .A1(n6762), .A2(n6761), .ZN(n10917) );
  AND2_X1 U5229 ( .A1(n6377), .A2(n9327), .ZN(n6386) );
  AND2_X1 U5230 ( .A1(n7917), .A2(n7202), .ZN(n7759) );
  NOR2_X1 U5231 ( .A1(n9361), .A2(n7749), .ZN(n9330) );
  OAI21_X1 U5232 ( .B1(n5983), .B2(n6174), .A(n5585), .ZN(n6178) );
  AND4_X1 U5233 ( .A1(n6712), .A2(n6711), .A3(n6710), .A4(n6709), .ZN(n8181)
         );
  NAND3_X2 U5234 ( .A1(n7732), .A2(n7731), .A3(n8235), .ZN(n7735) );
  AND4_X1 U5235 ( .A1(n6686), .A2(n6685), .A3(n6684), .A4(n6683), .ZN(n8015)
         );
  AOI21_X1 U5236 ( .B1(n5248), .B2(n5111), .A(n5144), .ZN(n5247) );
  AND4_X1 U5237 ( .A1(n6672), .A2(n6671), .A3(n6670), .A4(n6669), .ZN(n8798)
         );
  NAND4_X2 U5238 ( .A1(n6648), .A2(n6647), .A3(n6646), .A4(n6645), .ZN(n7077)
         );
  NAND2_X1 U5239 ( .A1(n5240), .A2(n5980), .ZN(n6160) );
  CLKBUF_X1 U5240 ( .A(n6853), .Z(n6951) );
  BUF_X2 U5241 ( .A(n5731), .Z(n6853) );
  NAND2_X1 U5242 ( .A1(n6667), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6648) );
  OR2_X1 U5243 ( .A1(n5092), .A2(n7360), .ZN(n6666) );
  INV_X2 U5244 ( .A(n6676), .ZN(n6890) );
  NAND3_X1 U5245 ( .A1(n6093), .A2(n6092), .A3(n6091), .ZN(n9405) );
  CLKBUF_X3 U5246 ( .A(n6667), .Z(n6898) );
  NAND4_X1 U5247 ( .A1(n6121), .A2(n6120), .A3(n6119), .A4(n6118), .ZN(n9402)
         );
  NAND4_X1 U5248 ( .A1(n6106), .A2(n6105), .A3(n6104), .A4(n6103), .ZN(n9403)
         );
  MUX2_X1 U5249 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10587), .S(n7410), .Z(n7976)
         );
  NAND2_X1 U5250 ( .A1(n7152), .A2(n7157), .ZN(n8653) );
  NAND2_X1 U5251 ( .A1(n10580), .A2(n6564), .ZN(n8790) );
  CLKBUF_X1 U5252 ( .A(n7150), .Z(n8788) );
  MUX2_X1 U5253 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6563), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n6564) );
  MUX2_X1 U5254 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7156), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n7157) );
  OR2_X1 U5255 ( .A1(n7479), .A2(n5477), .ZN(n5476) );
  AOI21_X1 U5256 ( .B1(n5984), .B2(n5586), .A(n5142), .ZN(n5585) );
  CLKBUF_X1 U5257 ( .A(n5957), .Z(n9256) );
  CLKBUF_X1 U5258 ( .A(n5956), .Z(n5959) );
  XNOR2_X1 U5259 ( .A(n6990), .B(n6543), .ZN(n7525) );
  NAND2_X1 U5260 ( .A1(n10580), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6561) );
  XNOR2_X1 U5261 ( .A(n5952), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5956) );
  NOR2_X1 U5262 ( .A1(n5782), .A2(n5781), .ZN(n5783) );
  XNOR2_X1 U5263 ( .A(n6987), .B(P1_IR_REG_21__SCAN_IN), .ZN(n7161) );
  XNOR2_X1 U5264 ( .A(n5955), .B(n5954), .ZN(n5957) );
  OAI21_X1 U5265 ( .B1(n6137), .B2(n5345), .A(n6148), .ZN(n5580) );
  OAI21_X1 U5266 ( .B1(n5594), .B2(n6084), .A(n5969), .ZN(n6107) );
  INV_X1 U5267 ( .A(n6544), .ZN(n6554) );
  NAND2_X1 U5268 ( .A1(n5779), .A2(n5713), .ZN(n5784) );
  OR2_X1 U5269 ( .A1(n6225), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U5270 ( .A1(n5953), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U5271 ( .A1(n9781), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5952) );
  XNOR2_X1 U5272 ( .A(n5831), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10721) );
  NAND2_X1 U5273 ( .A1(n5346), .A2(SI_4_), .ZN(n5978) );
  XNOR2_X1 U5274 ( .A(n5346), .B(n8884), .ZN(n6137) );
  NAND2_X2 U5275 ( .A1(n7362), .A2(P1_U3086), .ZN(n8793) );
  AND2_X1 U5276 ( .A1(n5774), .A2(n5778), .ZN(n5775) );
  AND2_X1 U5277 ( .A1(n5705), .A2(n6543), .ZN(n5403) );
  NOR2_X1 U5278 ( .A1(n5750), .A2(n5670), .ZN(n5669) );
  AND2_X1 U5279 ( .A1(n5765), .A2(n5764), .ZN(n5774) );
  AND2_X1 U5280 ( .A1(n6553), .A2(n5706), .ZN(n5705) );
  OAI21_X1 U5281 ( .B1(P1_RD_REG_SCAN_IN), .B2(P2_ADDR_REG_19__SCAN_IN), .A(
        n5596), .ZN(n5595) );
  AND2_X1 U5282 ( .A1(n5733), .A2(n5732), .ZN(n5807) );
  NAND4_X1 U5283 ( .A1(n5505), .A2(n5504), .A3(n5503), .A4(n5502), .ZN(n6535)
         );
  NOR2_X2 U5284 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5799) );
  INV_X1 U5285 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5596) );
  INV_X4 U5286 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5287 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6541) );
  INV_X1 U5288 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5803) );
  NOR2_X1 U5289 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5732) );
  NOR2_X1 U5290 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5733) );
  INV_X1 U5291 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9211) );
  INV_X1 U5292 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9212) );
  NOR2_X1 U5293 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5505) );
  NOR2_X1 U5294 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5389) );
  OR2_X1 U5295 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5813) );
  INV_X1 U5296 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9221) );
  INV_X1 U5297 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5747) );
  NOR2_X1 U5298 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n5562) );
  AOI21_X2 U5299 ( .B1(n8636), .B2(n8635), .A(n8634), .ZN(n10254) );
  NAND2_X1 U5300 ( .A1(n5783), .A2(n5784), .ZN(n5087) );
  NAND2_X1 U5301 ( .A1(n5783), .A2(n5784), .ZN(n5088) );
  NAND2_X1 U5302 ( .A1(n5783), .A2(n5784), .ZN(n5191) );
  AND2_X1 U5303 ( .A1(n7213), .A2(n7191), .ZN(n5487) );
  NAND2_X1 U5304 ( .A1(n7634), .A2(n7633), .ZN(n6450) );
  AND2_X1 U5305 ( .A1(n6574), .A2(n8790), .ZN(n6668) );
  NOR2_X2 U5306 ( .A1(n6236), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6249) );
  NAND2_X1 U5307 ( .A1(n7151), .A2(n7150), .ZN(n5089) );
  NAND2_X1 U5308 ( .A1(n7151), .A2(n7150), .ZN(n5090) );
  NAND2_X4 U5309 ( .A1(n7511), .A2(n7513), .ZN(n7808) );
  NAND2_X4 U5310 ( .A1(n7495), .A2(n7160), .ZN(n7511) );
  NOR2_X2 U5311 ( .A1(n6261), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6273) );
  NOR2_X2 U5312 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(n6363), .ZN(n6377) );
  NAND2_X1 U5313 ( .A1(n5090), .A2(n7362), .ZN(n5092) );
  INV_X1 U5314 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5761) );
  OR2_X1 U5315 ( .A1(n8811), .A2(n9316), .ZN(n7264) );
  OR2_X1 U5316 ( .A1(n9312), .A2(n8806), .ZN(n7252) );
  NAND2_X1 U5317 ( .A1(n6436), .A2(n6435), .ZN(n6548) );
  INV_X1 U5318 ( .A(n5542), .ZN(n5541) );
  INV_X1 U5319 ( .A(n7262), .ZN(n7256) );
  NAND2_X1 U5320 ( .A1(n5298), .A2(n5297), .ZN(n5296) );
  AND2_X1 U5321 ( .A1(n7328), .A2(n7320), .ZN(n7350) );
  NOR2_X1 U5322 ( .A1(n5547), .A2(n6317), .ZN(n5546) );
  INV_X1 U5323 ( .A(n5549), .ZN(n5547) );
  INV_X1 U5324 ( .A(n6267), .ZN(n6015) );
  NAND2_X1 U5325 ( .A1(n6000), .A2(n5999), .ZN(n6003) );
  INV_X1 U5326 ( .A(n5957), .ZN(n5958) );
  XNOR2_X1 U5327 ( .A(n5571), .B(n7371), .ZN(n10697) );
  OR2_X1 U5328 ( .A1(n6510), .A2(n9550), .ZN(n7303) );
  OR2_X1 U5329 ( .A1(n9657), .A2(n9636), .ZN(n7268) );
  OR2_X1 U5330 ( .A1(n9674), .A2(n9655), .ZN(n7265) );
  OR2_X1 U5331 ( .A1(n8111), .A2(n8449), .ZN(n7218) );
  INV_X1 U5332 ( .A(n5791), .ZN(n5668) );
  INV_X1 U5333 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U5334 ( .A1(n5743), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6446) );
  INV_X1 U5335 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5734) );
  AND2_X1 U5336 ( .A1(n7544), .A2(n7512), .ZN(n7510) );
  NAND2_X1 U5337 ( .A1(n5451), .A2(n7974), .ZN(n5456) );
  NAND2_X1 U5338 ( .A1(n5453), .A2(n5452), .ZN(n5451) );
  OR2_X1 U5339 ( .A1(n10491), .A2(n5413), .ZN(n5412) );
  OR2_X1 U5340 ( .A1(n10514), .A2(n9986), .ZN(n10239) );
  OR2_X1 U5341 ( .A1(n7507), .A2(n7512), .ZN(n7974) );
  NAND2_X1 U5342 ( .A1(n6415), .A2(n6414), .ZN(n6432) );
  NAND2_X1 U5343 ( .A1(n5258), .A2(n5257), .ZN(n6399) );
  AOI21_X1 U5344 ( .B1(n5107), .B2(n5263), .A(n5183), .ZN(n5257) );
  NOR2_X1 U5345 ( .A1(n6030), .A2(n5593), .ZN(n5592) );
  INV_X1 U5346 ( .A(n6025), .ZN(n5593) );
  NAND2_X1 U5347 ( .A1(n5608), .A2(n5103), .ZN(n6021) );
  INV_X1 U5348 ( .A(n6282), .ZN(n5607) );
  AND2_X1 U5349 ( .A1(n6025), .A2(n6024), .ZN(n6295) );
  NAND2_X1 U5350 ( .A1(n5994), .A2(n5993), .ZN(n6207) );
  NAND2_X1 U5351 ( .A1(n9345), .A2(n8823), .ZN(n8824) );
  OAI21_X1 U5352 ( .B1(n9280), .B2(n5121), .A(n5237), .ZN(n5236) );
  NAND2_X1 U5353 ( .A1(n9280), .A2(n5239), .ZN(n5237) );
  AND2_X1 U5354 ( .A1(n7730), .A2(n7354), .ZN(n7739) );
  AOI21_X1 U5355 ( .B1(n5632), .B2(n5634), .A(n5220), .ZN(n5219) );
  INV_X1 U5356 ( .A(n5632), .ZN(n5221) );
  INV_X1 U5357 ( .A(n8710), .ZN(n5220) );
  NAND2_X1 U5358 ( .A1(n5601), .A2(n5372), .ZN(n5278) );
  NAND2_X1 U5359 ( .A1(n7349), .A2(n5373), .ZN(n5372) );
  NAND2_X1 U5360 ( .A1(n5605), .A2(n6465), .ZN(n5601) );
  AND2_X1 U5361 ( .A1(n7328), .A2(n5186), .ZN(n5373) );
  NAND2_X1 U5362 ( .A1(n5600), .A2(n5124), .ZN(n5599) );
  INV_X1 U5363 ( .A(n5602), .ZN(n5600) );
  XNOR2_X1 U5364 ( .A(n5875), .B(n10702), .ZN(n10694) );
  INV_X1 U5365 ( .A(n5571), .ZN(n5823) );
  OR2_X1 U5366 ( .A1(n7857), .A2(n10716), .ZN(n5483) );
  NAND2_X1 U5367 ( .A1(n5878), .A2(n5481), .ZN(n5480) );
  INV_X1 U5368 ( .A(n7857), .ZN(n5481) );
  NOR2_X1 U5369 ( .A1(n7845), .A2(n5836), .ZN(n5837) );
  AND2_X1 U5370 ( .A1(n7392), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U5371 ( .A1(n5862), .A2(n5860), .ZN(n5564) );
  XNOR2_X1 U5372 ( .A(n5098), .B(n6297), .ZN(n9497) );
  AOI22_X1 U5373 ( .A1(n9621), .A2(n6370), .B1(n9611), .B2(n9714), .ZN(n9610)
         );
  INV_X1 U5374 ( .A(n5349), .ZN(n5348) );
  NAND2_X1 U5375 ( .A1(n8724), .A2(n6459), .ZN(n5350) );
  OAI21_X1 U5376 ( .B1(n6458), .B2(n5351), .A(n7264), .ZN(n5349) );
  AND4_X1 U5377 ( .A1(n6279), .A2(n6278), .A3(n6277), .A4(n6276), .ZN(n9307)
         );
  OAI21_X1 U5378 ( .B1(n8088), .B2(n5556), .A(n5203), .ZN(n6243) );
  AOI21_X1 U5379 ( .B1(n5204), .B2(n5555), .A(n6454), .ZN(n5203) );
  NAND2_X1 U5380 ( .A1(n8268), .A2(n7240), .ZN(n5365) );
  NAND2_X1 U5381 ( .A1(n5769), .A2(n5768), .ZN(n7722) );
  AND2_X1 U5382 ( .A1(n5767), .A2(n6488), .ZN(n5768) );
  NAND2_X1 U5383 ( .A1(n5215), .A2(n5113), .ZN(n5861) );
  AND2_X1 U5384 ( .A1(n7809), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7358) );
  NAND2_X1 U5385 ( .A1(n6558), .A2(n6557), .ZN(n10226) );
  OR2_X1 U5386 ( .A1(n10396), .A2(n10263), .ZN(n5719) );
  NAND2_X1 U5387 ( .A1(n7107), .A2(n5530), .ZN(n5529) );
  NAND2_X1 U5388 ( .A1(n7022), .A2(n7104), .ZN(n5530) );
  INV_X1 U5389 ( .A(n7410), .ZN(n6894) );
  NAND2_X1 U5390 ( .A1(n5089), .A2(n5417), .ZN(n6676) );
  NAND2_X1 U5391 ( .A1(n5090), .A2(n7362), .ZN(n6692) );
  AND2_X1 U5392 ( .A1(n7511), .A2(n7358), .ZN(n10573) );
  XNOR2_X1 U5393 ( .A(n6432), .B(n6431), .ZN(n8787) );
  AND2_X1 U5394 ( .A1(n5705), .A2(n5400), .ZN(n5401) );
  AND2_X1 U5395 ( .A1(n6543), .A2(n5402), .ZN(n5400) );
  INV_X1 U5396 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U5397 ( .A1(n5212), .A2(n5131), .ZN(n9271) );
  NAND2_X1 U5398 ( .A1(n9306), .A2(n5622), .ZN(n5212) );
  NOR2_X1 U5399 ( .A1(n5564), .A2(n9501), .ZN(n9511) );
  INV_X1 U5400 ( .A(n9748), .ZN(n9555) );
  AOI21_X1 U5401 ( .B1(n6821), .B2(n6820), .A(n6819), .ZN(n6863) );
  AND2_X1 U5402 ( .A1(n7024), .A2(n7107), .ZN(n5327) );
  NAND2_X1 U5403 ( .A1(n5336), .A2(n10237), .ZN(n5335) );
  NAND2_X1 U5404 ( .A1(n6921), .A2(n6920), .ZN(n5336) );
  OR2_X1 U5405 ( .A1(n6935), .A2(n6993), .ZN(n6923) );
  NAND2_X1 U5406 ( .A1(n10242), .A2(n7547), .ZN(n5340) );
  INV_X1 U5407 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9169) );
  INV_X1 U5408 ( .A(n7270), .ZN(n5319) );
  NOR2_X1 U5409 ( .A1(n7348), .A2(n7347), .ZN(n5286) );
  INV_X1 U5410 ( .A(n7349), .ZN(n5285) );
  NOR2_X1 U5411 ( .A1(n5366), .A2(n5367), .ZN(n5364) );
  INV_X1 U5412 ( .A(n7240), .ZN(n5367) );
  INV_X1 U5413 ( .A(n8740), .ZN(n5255) );
  AND2_X1 U5414 ( .A1(n9802), .A2(n5711), .ZN(n5256) );
  INV_X1 U5415 ( .A(n5446), .ZN(n5252) );
  AOI21_X1 U5416 ( .B1(n9802), .B2(n8745), .A(n5136), .ZN(n5446) );
  INV_X1 U5417 ( .A(n5441), .ZN(n5440) );
  OAI21_X1 U5418 ( .B1(n8328), .B2(n5442), .A(n8565), .ZN(n5441) );
  INV_X1 U5419 ( .A(n8333), .ZN(n5442) );
  INV_X1 U5420 ( .A(SI_17_), .ZN(n9064) );
  INV_X1 U5421 ( .A(SI_14_), .ZN(n9069) );
  INV_X1 U5422 ( .A(SI_12_), .ZN(n8869) );
  INV_X1 U5423 ( .A(SI_10_), .ZN(n9078) );
  OAI211_X1 U5424 ( .C1(n8437), .C2(n5145), .A(n5223), .B(n5104), .ZN(n5222)
         );
  OR2_X1 U5425 ( .A1(n5712), .A2(n5224), .ZN(n5223) );
  NOR2_X1 U5426 ( .A1(n7327), .A2(n7326), .ZN(n7330) );
  INV_X1 U5427 ( .A(n5869), .ZN(n5471) );
  NOR2_X1 U5428 ( .A1(n7296), .A2(n5386), .ZN(n5385) );
  INV_X1 U5429 ( .A(n6462), .ZN(n5386) );
  NOR2_X1 U5430 ( .A1(n6396), .A2(n6395), .ZN(n9561) );
  AND2_X1 U5431 ( .A1(n9584), .A2(n9386), .ZN(n6395) );
  NOR2_X1 U5432 ( .A1(n9574), .A2(n5126), .ZN(n6396) );
  OR2_X1 U5433 ( .A1(n8760), .A2(n9307), .ZN(n7175) );
  AND2_X1 U5434 ( .A1(n5361), .A2(n8461), .ZN(n5368) );
  NAND2_X1 U5435 ( .A1(n8266), .A2(n7240), .ZN(n5361) );
  NAND2_X1 U5436 ( .A1(n5558), .A2(n6219), .ZN(n5557) );
  INV_X1 U5437 ( .A(n7337), .ZN(n5558) );
  NOR2_X1 U5438 ( .A1(n8101), .A2(n5560), .ZN(n5559) );
  INV_X1 U5439 ( .A(n6206), .ZN(n5560) );
  INV_X1 U5440 ( .A(n7200), .ZN(n5358) );
  INV_X1 U5441 ( .A(n7917), .ZN(n5357) );
  AND2_X1 U5442 ( .A1(n5761), .A2(n5760), .ZN(n5765) );
  NAND2_X1 U5443 ( .A1(n5742), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5786) );
  INV_X1 U5444 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5814) );
  INV_X1 U5445 ( .A(n5430), .ZN(n5429) );
  OAI21_X1 U5446 ( .B1(n5432), .B2(n5431), .A(n9972), .ZN(n5430) );
  NAND2_X1 U5447 ( .A1(n5455), .A2(n5456), .ZN(n5454) );
  INV_X1 U5448 ( .A(n7510), .ZN(n5455) );
  NAND2_X1 U5449 ( .A1(n10290), .A2(n5414), .ZN(n5413) );
  OR2_X1 U5450 ( .A1(n10506), .A2(n10305), .ZN(n7041) );
  NAND2_X1 U5451 ( .A1(n10362), .A2(n5515), .ZN(n5514) );
  INV_X1 U5452 ( .A(n10238), .ZN(n5515) );
  NOR2_X1 U5453 ( .A1(n10514), .A2(n5392), .ZN(n5391) );
  INV_X1 U5454 ( .A(n5393), .ZN(n5392) );
  NOR2_X1 U5455 ( .A1(n10520), .A2(n10525), .ZN(n5393) );
  OR2_X1 U5456 ( .A1(n10531), .A2(n10263), .ZN(n7044) );
  INV_X1 U5457 ( .A(n5690), .ZN(n5689) );
  OR2_X1 U5458 ( .A1(n10556), .A2(n10465), .ZN(n7018) );
  NOR2_X1 U5459 ( .A1(n5528), .A2(n8366), .ZN(n5672) );
  OR2_X1 U5460 ( .A1(n8619), .A2(n8746), .ZN(n10939) );
  AND2_X1 U5461 ( .A1(n5528), .A2(n7008), .ZN(n5527) );
  NOR2_X1 U5462 ( .A1(n5680), .A2(n8186), .ZN(n5677) );
  INV_X1 U5463 ( .A(n10890), .ZN(n5680) );
  OAI21_X1 U5464 ( .B1(n7088), .B2(n5536), .A(n7987), .ZN(n5532) );
  OR2_X1 U5465 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n6559) );
  INV_X1 U5466 ( .A(n6559), .ZN(n5702) );
  OAI21_X1 U5467 ( .B1(n6399), .B2(n6398), .A(n6397), .ZN(n6413) );
  NOR2_X1 U5468 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5706) );
  NAND2_X1 U5469 ( .A1(n6988), .A2(n6543), .ZN(n6544) );
  AND2_X1 U5470 ( .A1(n6055), .A2(n6054), .ZN(n6373) );
  NAND2_X1 U5471 ( .A1(n6544), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6987) );
  INV_X1 U5472 ( .A(n6318), .ZN(n5591) );
  XNOR2_X1 U5473 ( .A(n6013), .B(n6012), .ZN(n6267) );
  INV_X1 U5474 ( .A(n5997), .ZN(n5617) );
  INV_X1 U5475 ( .A(n5616), .ZN(n5615) );
  OAI21_X1 U5476 ( .B1(n6208), .B2(n5111), .A(n6003), .ZN(n5616) );
  INV_X1 U5477 ( .A(n6177), .ZN(n5584) );
  INV_X1 U5478 ( .A(n5655), .ZN(n5653) );
  NAND2_X1 U5479 ( .A1(n5659), .A2(n5167), .ZN(n5655) );
  AOI21_X1 U5480 ( .B1(n5635), .B2(n5633), .A(n8707), .ZN(n5632) );
  INV_X1 U5481 ( .A(n8663), .ZN(n5633) );
  AND2_X1 U5482 ( .A1(n7743), .A2(n7741), .ZN(n5666) );
  INV_X1 U5483 ( .A(n9304), .ZN(n5629) );
  NAND2_X1 U5484 ( .A1(n5664), .A2(n5665), .ZN(n5662) );
  NAND2_X1 U5485 ( .A1(n7764), .A2(n9402), .ZN(n5665) );
  OR2_X1 U5486 ( .A1(n8057), .A2(n8056), .ZN(n5214) );
  INV_X1 U5487 ( .A(n5381), .ZN(n5380) );
  AND2_X1 U5488 ( .A1(n5959), .A2(n9256), .ZN(n6115) );
  NOR2_X1 U5489 ( .A1(n7440), .A2(n7439), .ZN(n7438) );
  INV_X1 U5490 ( .A(n5819), .ZN(n5309) );
  OR2_X1 U5491 ( .A1(n10676), .A2(n7480), .ZN(n5477) );
  NAND2_X1 U5492 ( .A1(n5874), .A2(n5475), .ZN(n5474) );
  INV_X1 U5493 ( .A(n10676), .ZN(n5475) );
  NOR2_X1 U5494 ( .A1(n10697), .A2(n10698), .ZN(n10696) );
  NAND2_X1 U5495 ( .A1(n5293), .A2(n5291), .ZN(n7461) );
  OR2_X1 U5496 ( .A1(n10697), .A2(n5155), .ZN(n5293) );
  NAND2_X1 U5497 ( .A1(n5824), .A2(n5292), .ZN(n5291) );
  NOR2_X1 U5498 ( .A1(n7461), .A2(n5827), .ZN(n5828) );
  NOR2_X1 U5499 ( .A1(n7467), .A2(n5826), .ZN(n5827) );
  XNOR2_X1 U5500 ( .A(n5828), .B(n10721), .ZN(n10713) );
  XNOR2_X1 U5501 ( .A(n5880), .B(n6195), .ZN(n8137) );
  NAND2_X1 U5502 ( .A1(n8207), .A2(n5563), .ZN(n5304) );
  NAND2_X1 U5503 ( .A1(n5306), .A2(n5563), .ZN(n5305) );
  NAND2_X1 U5504 ( .A1(n7404), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5563) );
  XNOR2_X1 U5505 ( .A(n5846), .B(n9442), .ZN(n9424) );
  NAND2_X1 U5506 ( .A1(n5460), .A2(n5459), .ZN(n5458) );
  INV_X1 U5507 ( .A(n9479), .ZN(n5459) );
  NAND2_X1 U5508 ( .A1(n9556), .A2(n7292), .ZN(n5387) );
  XNOR2_X1 U5509 ( .A(n9561), .B(n9566), .ZN(n9562) );
  NAND2_X1 U5510 ( .A1(n6372), .A2(n6371), .ZN(n9599) );
  NAND2_X1 U5511 ( .A1(n9618), .A2(n9601), .ZN(n6371) );
  NOR2_X1 U5512 ( .A1(n7280), .A2(n7169), .ZN(n5360) );
  NAND2_X1 U5513 ( .A1(n5463), .A2(n5461), .ZN(n9642) );
  AOI21_X1 U5514 ( .B1(n5099), .B2(n5468), .A(n5462), .ZN(n5461) );
  INV_X1 U5515 ( .A(n7268), .ZN(n5462) );
  AOI21_X1 U5516 ( .B1(n5093), .B2(n9676), .A(n5137), .ZN(n5553) );
  NAND2_X1 U5517 ( .A1(n5195), .A2(n5093), .ZN(n5194) );
  AOI21_X1 U5518 ( .B1(n7265), .B2(n5467), .A(n5466), .ZN(n5465) );
  INV_X1 U5519 ( .A(n7260), .ZN(n5467) );
  INV_X1 U5520 ( .A(n5195), .ZN(n9665) );
  NAND2_X1 U5521 ( .A1(n9665), .A2(n6330), .ZN(n9663) );
  AOI21_X1 U5522 ( .B1(n8725), .B2(n5550), .A(n5130), .ZN(n5549) );
  INV_X1 U5523 ( .A(n6293), .ZN(n5550) );
  AND2_X1 U5524 ( .A1(n7264), .A2(n7260), .ZN(n8699) );
  INV_X1 U5525 ( .A(n8724), .ZN(n5352) );
  AND4_X1 U5526 ( .A1(n6306), .A2(n6305), .A3(n6304), .A4(n6303), .ZN(n8809)
         );
  AND4_X1 U5527 ( .A1(n6292), .A2(n6291), .A3(n6290), .A4(n6289), .ZN(n8806)
         );
  AOI21_X1 U5528 ( .B1(n6266), .B2(n8461), .A(n5139), .ZN(n5542) );
  AND4_X1 U5529 ( .A1(n6265), .A2(n6264), .A3(n6263), .A4(n6262), .ZN(n8767)
         );
  INV_X1 U5530 ( .A(n8458), .ZN(n5543) );
  NAND2_X1 U5531 ( .A1(n7222), .A2(n6452), .ZN(n7237) );
  AND4_X1 U5532 ( .A1(n6254), .A2(n6253), .A3(n6252), .A4(n6251), .ZN(n8713)
         );
  INV_X1 U5533 ( .A(n9395), .ZN(n8473) );
  NOR2_X1 U5534 ( .A1(n5557), .A2(n8086), .ZN(n5205) );
  INV_X1 U5535 ( .A(n9394), .ZN(n8660) );
  NAND2_X1 U5536 ( .A1(n6199), .A2(n8114), .ZN(n6212) );
  AND2_X1 U5537 ( .A1(n8318), .A2(n8320), .ZN(n8101) );
  NAND2_X1 U5538 ( .A1(n8087), .A2(n5559), .ZN(n8096) );
  NAND2_X1 U5539 ( .A1(n6193), .A2(n6192), .ZN(n8088) );
  NAND2_X1 U5540 ( .A1(n8446), .A2(n6188), .ZN(n6193) );
  NAND2_X1 U5541 ( .A1(n8088), .A2(n6205), .ZN(n8087) );
  AND2_X1 U5542 ( .A1(n7915), .A2(n7203), .ZN(n7883) );
  AND2_X1 U5543 ( .A1(n7203), .A2(n7201), .ZN(n7920) );
  AOI22_X1 U5544 ( .A1(n6450), .A2(n5487), .B1(n7213), .B2(n5486), .ZN(n7681)
         );
  OR2_X1 U5545 ( .A1(n7749), .A2(n7306), .ZN(n9635) );
  INV_X1 U5546 ( .A(n7636), .ZN(n7633) );
  AND2_X1 U5547 ( .A1(n5637), .A2(n6489), .ZN(n8235) );
  NAND2_X1 U5548 ( .A1(n6487), .A2(n5127), .ZN(n5637) );
  NAND2_X1 U5549 ( .A1(n7749), .A2(n7739), .ZN(n9637) );
  NAND2_X1 U5550 ( .A1(n7311), .A2(n7310), .ZN(n7328) );
  NAND2_X1 U5551 ( .A1(n6438), .A2(n6437), .ZN(n6510) );
  NAND2_X1 U5552 ( .A1(n6310), .A2(n6309), .ZN(n8811) );
  AND2_X1 U5553 ( .A1(n6234), .A2(n6233), .ZN(n8471) );
  INV_X1 U5554 ( .A(n8726), .ZN(n9720) );
  INV_X1 U5555 ( .A(n7301), .ZN(n6321) );
  INV_X1 U5556 ( .A(n6475), .ZN(n6320) );
  NAND2_X1 U5557 ( .A1(n5754), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5759) );
  INV_X1 U5558 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5758) );
  INV_X1 U5559 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5735) );
  INV_X1 U5560 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5736) );
  XNOR2_X1 U5561 ( .A(n5805), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10702) );
  NAND2_X1 U5562 ( .A1(n5242), .A2(n10047), .ZN(n9930) );
  NAND2_X1 U5563 ( .A1(n8575), .A2(n8574), .ZN(n8603) );
  INV_X1 U5564 ( .A(n9984), .ZN(n5281) );
  INV_X1 U5565 ( .A(n9958), .ZN(n9959) );
  INV_X1 U5566 ( .A(n5456), .ZN(n5450) );
  NAND2_X1 U5567 ( .A1(n7507), .A2(n7525), .ZN(n7508) );
  AND4_X1 U5568 ( .A1(n6598), .A2(n6597), .A3(n6596), .A4(n6595), .ZN(n9986)
         );
  AND4_X1 U5569 ( .A1(n6736), .A2(n6735), .A3(n6734), .A4(n6733), .ZN(n8303)
         );
  NOR2_X1 U5570 ( .A1(n7872), .A2(n5171), .ZN(n7874) );
  INV_X1 U5571 ( .A(n10129), .ZN(n10124) );
  AND2_X1 U5572 ( .A1(n7039), .A2(n7125), .ZN(n10273) );
  OAI21_X1 U5573 ( .B1(n10303), .B2(n5519), .A(n5517), .ZN(n5523) );
  AOI21_X1 U5574 ( .B1(n5520), .B2(n10246), .A(n5518), .ZN(n5517) );
  INV_X1 U5575 ( .A(n5520), .ZN(n5519) );
  INV_X1 U5576 ( .A(n10247), .ZN(n5518) );
  OR2_X1 U5577 ( .A1(n10326), .A2(n10305), .ZN(n5722) );
  NAND2_X1 U5578 ( .A1(n10313), .A2(n5684), .ZN(n10298) );
  NOR2_X1 U5579 ( .A1(n5522), .A2(n5685), .ZN(n5684) );
  INV_X1 U5580 ( .A(n5722), .ZN(n5685) );
  OR2_X1 U5581 ( .A1(n10265), .A2(n10267), .ZN(n5721) );
  NAND2_X1 U5582 ( .A1(n10356), .A2(n10266), .ZN(n10268) );
  NAND2_X1 U5583 ( .A1(n10421), .A2(n5697), .ZN(n5696) );
  NOR2_X1 U5584 ( .A1(n10410), .A2(n5698), .ZN(n5697) );
  NOR2_X1 U5585 ( .A1(n10403), .A2(n10531), .ZN(n10393) );
  AND2_X1 U5586 ( .A1(n7045), .A2(n10236), .ZN(n10410) );
  OR2_X1 U5587 ( .A1(n11032), .A2(n10433), .ZN(n5718) );
  AND2_X1 U5588 ( .A1(n10543), .A2(n10258), .ZN(n10259) );
  AND4_X1 U5589 ( .A1(n6875), .A2(n6874), .A3(n6873), .A4(n6872), .ZN(n10450)
         );
  NAND2_X1 U5590 ( .A1(n5531), .A2(n7021), .ZN(n10461) );
  INV_X1 U5591 ( .A(n10459), .ZN(n5531) );
  NOR2_X1 U5592 ( .A1(n10556), .A2(n5693), .ZN(n5692) );
  NAND2_X1 U5593 ( .A1(n10469), .A2(n5691), .ZN(n5690) );
  INV_X1 U5594 ( .A(n5692), .ZN(n5691) );
  NOR2_X1 U5595 ( .A1(n10547), .A2(n10548), .ZN(n10546) );
  AOI21_X1 U5596 ( .B1(n7058), .B2(n5511), .A(n5510), .ZN(n5509) );
  INV_X1 U5597 ( .A(n7015), .ZN(n5511) );
  INV_X1 U5598 ( .A(n7057), .ZN(n5510) );
  INV_X1 U5599 ( .A(n10462), .ZN(n10552) );
  NOR2_X1 U5600 ( .A1(n10948), .A2(n9799), .ZN(n8644) );
  OR2_X1 U5601 ( .A1(n10957), .A2(n10094), .ZN(n8548) );
  NAND2_X1 U5602 ( .A1(n8427), .A2(n8583), .ZN(n7008) );
  NAND2_X1 U5603 ( .A1(n7009), .A2(n5527), .ZN(n10943) );
  NOR2_X1 U5604 ( .A1(n7536), .A2(n7535), .ZN(n7948) );
  OR2_X1 U5605 ( .A1(n5092), .A2(n7385), .ZN(n6678) );
  AND2_X1 U5606 ( .A1(n7542), .A2(n7541), .ZN(n10941) );
  INV_X1 U5607 ( .A(n10219), .ZN(n7950) );
  NAND2_X1 U5608 ( .A1(n8788), .A2(n7656), .ZN(n10462) );
  NAND2_X1 U5609 ( .A1(n6572), .A2(n6571), .ZN(n10491) );
  AND2_X1 U5610 ( .A1(n7508), .A2(n7540), .ZN(n10557) );
  AND3_X1 U5611 ( .A1(n6708), .A2(n6707), .A3(n6706), .ZN(n10858) );
  NAND2_X1 U5612 ( .A1(n6704), .A2(n6890), .ZN(n6708) );
  NAND2_X1 U5613 ( .A1(n7410), .A2(n5416), .ZN(n5415) );
  OAI22_X1 U5614 ( .A1(n5115), .A2(n7362), .B1(n7377), .B2(n5417), .ZN(n5416)
         );
  INV_X1 U5615 ( .A(n10941), .ZN(n10821) );
  NAND2_X1 U5616 ( .A1(n6548), .A2(n5268), .ZN(n5267) );
  NOR2_X1 U5617 ( .A1(n6978), .A2(n5270), .ZN(n5268) );
  AOI21_X1 U5618 ( .B1(n5266), .B2(n5184), .A(n5265), .ZN(n5264) );
  INV_X1 U5619 ( .A(n6977), .ZN(n5265) );
  INV_X1 U5620 ( .A(n6978), .ZN(n5266) );
  XNOR2_X1 U5621 ( .A(n6979), .B(n6978), .ZN(n9258) );
  AOI21_X1 U5622 ( .B1(n6548), .B2(n5269), .A(n5184), .ZN(n6979) );
  AND2_X1 U5623 ( .A1(n7154), .A2(n5404), .ZN(n7495) );
  NAND2_X1 U5624 ( .A1(n6064), .A2(n6050), .ZN(n6067) );
  XNOR2_X1 U5625 ( .A(n7147), .B(n9226), .ZN(n7809) );
  NAND2_X1 U5626 ( .A1(n6333), .A2(n6332), .ZN(n6335) );
  NAND2_X1 U5627 ( .A1(n5587), .A2(n6029), .ZN(n6319) );
  NAND2_X1 U5628 ( .A1(n6026), .A2(n5592), .ZN(n5587) );
  NAND2_X1 U5629 ( .A1(n5608), .A2(n5609), .ZN(n6283) );
  OR2_X1 U5630 ( .A1(n6740), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6808) );
  XNOR2_X1 U5631 ( .A(n6705), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7706) );
  XNOR2_X1 U5632 ( .A(n6173), .B(n6174), .ZN(n6704) );
  NAND2_X1 U5633 ( .A1(n5983), .A2(n5982), .ZN(n6173) );
  NOR2_X1 U5634 ( .A1(n5300), .A2(n7297), .ZN(n5299) );
  NAND2_X2 U5635 ( .A1(n5087), .A2(n5864), .ZN(n6475) );
  AND4_X1 U5636 ( .A1(n6369), .A2(n6368), .A3(n6367), .A4(n6366), .ZN(n9638)
         );
  AND4_X1 U5637 ( .A1(n6218), .A2(n6217), .A3(n6216), .A4(n6215), .ZN(n8325)
         );
  NOR2_X1 U5638 ( .A1(n5102), .A2(n9355), .ZN(n5232) );
  INV_X1 U5639 ( .A(n5239), .ZN(n5235) );
  NAND2_X1 U5640 ( .A1(n5236), .A2(n5238), .ZN(n5234) );
  NAND2_X1 U5641 ( .A1(n9280), .A2(n9279), .ZN(n5238) );
  NAND2_X1 U5642 ( .A1(n5618), .A2(n6385), .ZN(n6393) );
  NAND2_X1 U5643 ( .A1(n8632), .A2(n7308), .ZN(n5618) );
  NAND2_X1 U5644 ( .A1(n8805), .A2(n5720), .ZN(n9306) );
  OR2_X1 U5645 ( .A1(n8804), .A2(n9307), .ZN(n5720) );
  INV_X1 U5646 ( .A(n9764), .ZN(n9334) );
  NAND2_X1 U5647 ( .A1(n8113), .A2(n8112), .ZN(n8254) );
  AND4_X1 U5648 ( .A1(n6329), .A2(n6328), .A3(n6327), .A4(n6326), .ZN(n9655)
         );
  INV_X1 U5649 ( .A(n9588), .ZN(n9612) );
  NOR2_X1 U5650 ( .A1(n5828), .A2(n10721), .ZN(n5829) );
  NOR2_X1 U5651 ( .A1(n10713), .A2(n10876), .ZN(n10712) );
  AND2_X1 U5652 ( .A1(n5485), .A2(n5484), .ZN(n7858) );
  NAND2_X1 U5653 ( .A1(n5482), .A2(n5480), .ZN(n7856) );
  OAI21_X1 U5654 ( .B1(n10713), .B2(n5569), .A(n5310), .ZN(n7845) );
  OR2_X1 U5655 ( .A1(n7846), .A2(n10876), .ZN(n5569) );
  NAND2_X1 U5656 ( .A1(n5829), .A2(n5570), .ZN(n5310) );
  INV_X1 U5657 ( .A(n7846), .ZN(n5570) );
  INV_X1 U5658 ( .A(n5495), .ZN(n9436) );
  NAND2_X1 U5659 ( .A1(n9507), .A2(n10729), .ZN(n5577) );
  AOI21_X1 U5660 ( .B1(n9505), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n5579), .ZN(
        n5578) );
  NOR2_X1 U5661 ( .A1(n9521), .A2(n9506), .ZN(n5579) );
  AOI21_X1 U5662 ( .B1(n9528), .B2(n9527), .A(n9526), .ZN(n9529) );
  NOR2_X1 U5663 ( .A1(n9496), .A2(n5892), .ZN(n9510) );
  INV_X1 U5664 ( .A(n10734), .ZN(n9505) );
  NAND2_X1 U5665 ( .A1(n9509), .A2(n5893), .ZN(n5498) );
  OAI22_X1 U5666 ( .A1(n5862), .A2(n5289), .B1(n8701), .B2(n9527), .ZN(n5290)
         );
  NOR2_X1 U5667 ( .A1(n9522), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U5668 ( .A1(n7425), .A2(n5088), .ZN(n10717) );
  NAND2_X1 U5669 ( .A1(n6479), .A2(n9664), .ZN(n5207) );
  AOI21_X1 U5670 ( .B1(n9545), .B2(n8292), .A(n6478), .ZN(n5206) );
  INV_X1 U5671 ( .A(n9756), .ZN(n9584) );
  NAND2_X1 U5672 ( .A1(n9735), .A2(n9720), .ZN(n9738) );
  AND2_X1 U5673 ( .A1(n6418), .A2(n6417), .ZN(n9748) );
  AND2_X1 U5674 ( .A1(n6492), .A2(n6491), .ZN(n8238) );
  XNOR2_X1 U5675 ( .A(n5834), .B(n5833), .ZN(n7392) );
  NAND2_X1 U5676 ( .A1(n6897), .A2(n6896), .ZN(n10260) );
  INV_X1 U5677 ( .A(n10081), .ZN(n10064) );
  NAND2_X1 U5678 ( .A1(n7527), .A2(n10472), .ZN(n10073) );
  AOI21_X1 U5679 ( .B1(n7309), .B2(n6890), .A(n6982), .ZN(n10484) );
  OR2_X1 U5680 ( .A1(n6546), .A2(n9009), .ZN(n5287) );
  NAND2_X1 U5681 ( .A1(n5332), .A2(n5123), .ZN(n5331) );
  NAND2_X1 U5682 ( .A1(n6861), .A2(n7058), .ZN(n5332) );
  NAND2_X1 U5683 ( .A1(n6866), .A2(n7547), .ZN(n5330) );
  AOI21_X1 U5684 ( .B1(n6865), .B2(n7057), .A(n6864), .ZN(n6866) );
  INV_X1 U5685 ( .A(n6889), .ZN(n5329) );
  NAND2_X1 U5686 ( .A1(n7222), .A2(n5314), .ZN(n5313) );
  NAND2_X1 U5687 ( .A1(n7238), .A2(n7306), .ZN(n5316) );
  NAND2_X1 U5688 ( .A1(n6916), .A2(n6915), .ZN(n6921) );
  MUX2_X1 U5689 ( .A(n6914), .B(n6913), .S(n7547), .Z(n6915) );
  NAND2_X1 U5690 ( .A1(n5337), .A2(n5333), .ZN(n6935) );
  NAND2_X1 U5691 ( .A1(n5335), .A2(n5334), .ZN(n5333) );
  AND2_X1 U5692 ( .A1(n7043), .A2(n7547), .ZN(n5334) );
  NAND2_X1 U5693 ( .A1(n5311), .A2(n7254), .ZN(n7262) );
  NOR2_X1 U5694 ( .A1(n5466), .A2(n5322), .ZN(n5321) );
  NAND2_X1 U5695 ( .A1(n7260), .A2(n7306), .ZN(n5322) );
  AND2_X1 U5696 ( .A1(n7264), .A2(n7739), .ZN(n5324) );
  NAND2_X1 U5697 ( .A1(n5299), .A2(n7299), .ZN(n5298) );
  INV_X1 U5698 ( .A(n7298), .ZN(n5297) );
  OAI21_X1 U5699 ( .B1(n5341), .B2(n5339), .A(n7040), .ZN(n5338) );
  AOI21_X1 U5700 ( .B1(n6937), .B2(n6997), .A(n5340), .ZN(n5339) );
  INV_X1 U5701 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9168) );
  INV_X1 U5702 ( .A(SI_9_), .ZN(n9077) );
  INV_X1 U5703 ( .A(n8469), .ZN(n5224) );
  NOR2_X1 U5704 ( .A1(n10480), .A2(n5398), .ZN(n5397) );
  INV_X1 U5705 ( .A(n5399), .ZN(n5398) );
  NOR2_X1 U5706 ( .A1(n8583), .A2(n8345), .ZN(n5409) );
  INV_X1 U5707 ( .A(SI_21_), .ZN(n9059) );
  NAND2_X1 U5708 ( .A1(n6017), .A2(n6016), .ZN(n6020) );
  NAND2_X1 U5709 ( .A1(n6207), .A2(n5247), .ZN(n5245) );
  NAND2_X1 U5710 ( .A1(n5598), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U5711 ( .A1(n5318), .A2(n5317), .ZN(n7274) );
  AND2_X1 U5712 ( .A1(n9641), .A2(n7269), .ZN(n5317) );
  OR2_X1 U5713 ( .A1(n6393), .A2(n9602), .ZN(n7285) );
  OR2_X1 U5714 ( .A1(n5628), .A2(n5717), .ZN(n5626) );
  AND2_X1 U5715 ( .A1(n9315), .A2(n5629), .ZN(n5628) );
  OAI21_X1 U5716 ( .B1(n7348), .B2(n5382), .A(n7322), .ZN(n5381) );
  NAND2_X1 U5717 ( .A1(n5387), .A2(n6463), .ZN(n5382) );
  NOR2_X1 U5718 ( .A1(n5383), .A2(n5378), .ZN(n5377) );
  INV_X1 U5719 ( .A(n5385), .ZN(n5378) );
  NAND2_X1 U5720 ( .A1(n5384), .A2(n6463), .ZN(n5383) );
  NAND2_X1 U5721 ( .A1(n5606), .A2(n7351), .ZN(n5605) );
  NAND2_X1 U5722 ( .A1(n5284), .A2(n8122), .ZN(n5606) );
  AOI21_X1 U5723 ( .B1(n5604), .B2(n5603), .A(n7319), .ZN(n5602) );
  OR2_X1 U5724 ( .A1(n7350), .A2(n7349), .ZN(n7319) );
  NOR2_X1 U5725 ( .A1(n7438), .A2(n5872), .ZN(n5873) );
  AND2_X1 U5726 ( .A1(n7363), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5872) );
  OR2_X1 U5727 ( .A1(n10678), .A2(n5157), .ZN(n5571) );
  INV_X1 U5728 ( .A(n7462), .ZN(n5292) );
  INV_X1 U5729 ( .A(n5838), .ZN(n5306) );
  OR2_X1 U5730 ( .A1(n9334), .A2(n9588), .ZN(n7279) );
  OR2_X1 U5731 ( .A1(n9719), .A2(n9654), .ZN(n7271) );
  NAND2_X1 U5732 ( .A1(n5544), .A2(n5545), .ZN(n5195) );
  AOI21_X1 U5733 ( .B1(n5546), .B2(n6458), .A(n5134), .ZN(n5545) );
  OR2_X1 U5734 ( .A1(n6324), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6338) );
  AOI21_X1 U5735 ( .B1(n5542), .B2(n5540), .A(n5539), .ZN(n5538) );
  INV_X1 U5736 ( .A(n8626), .ZN(n5539) );
  INV_X1 U5737 ( .A(n6266), .ZN(n5540) );
  OR2_X1 U5738 ( .A1(n5368), .A2(n5366), .ZN(n5362) );
  INV_X1 U5739 ( .A(n5205), .ZN(n5204) );
  NAND2_X1 U5740 ( .A1(n7234), .A2(n8318), .ZN(n7222) );
  AND2_X1 U5741 ( .A1(n5159), .A2(n6127), .ZN(n5200) );
  AND2_X1 U5742 ( .A1(n5775), .A2(n5951), .ZN(n5561) );
  NAND2_X1 U5743 ( .A1(n5776), .A2(n5775), .ZN(n5780) );
  INV_X1 U5744 ( .A(n5780), .ZN(n5782) );
  NAND2_X1 U5745 ( .A1(n5753), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5771) );
  INV_X1 U5746 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U5747 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), 
        .ZN(n5216) );
  OR2_X1 U5748 ( .A1(n5749), .A2(n5806), .ZN(n5740) );
  NAND2_X1 U5749 ( .A1(n5751), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5215) );
  NAND2_X1 U5750 ( .A1(n5253), .A2(n5251), .ZN(n9811) );
  NOR2_X1 U5751 ( .A1(n5133), .A2(n5252), .ZN(n5251) );
  AOI21_X1 U5752 ( .B1(n5440), .B2(n5442), .A(n5146), .ZN(n5438) );
  OR2_X1 U5753 ( .A1(n10776), .A2(n9860), .ZN(n7649) );
  INV_X1 U5754 ( .A(n9860), .ZN(n9948) );
  OR2_X1 U5755 ( .A1(n10491), .A2(n9960), .ZN(n7039) );
  NOR2_X1 U5756 ( .A1(n5521), .A2(n10291), .ZN(n5520) );
  NOR2_X1 U5757 ( .A1(n5522), .A2(n10246), .ZN(n5521) );
  OR2_X1 U5758 ( .A1(n10501), .A2(n10319), .ZN(n6992) );
  NAND2_X1 U5759 ( .A1(n6618), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6628) );
  AND2_X1 U5760 ( .A1(n6902), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6637) );
  NOR2_X1 U5761 ( .A1(n6900), .A2(n6899), .ZN(n6902) );
  NOR2_X1 U5762 ( .A1(n10556), .A2(n10255), .ZN(n5399) );
  NOR2_X1 U5763 ( .A1(n6855), .A2(n6854), .ZN(n6870) );
  NAND2_X1 U5764 ( .A1(n10927), .A2(n5409), .ZN(n5408) );
  INV_X1 U5765 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6772) );
  NAND2_X1 U5766 ( .A1(n7812), .A2(n7799), .ZN(n6679) );
  AND2_X1 U5767 ( .A1(n8644), .A2(n5395), .ZN(n10452) );
  AND2_X1 U5768 ( .A1(n5397), .A2(n5396), .ZN(n5395) );
  NAND2_X1 U5769 ( .A1(n8644), .A2(n5397), .ZN(n10476) );
  NOR2_X1 U5770 ( .A1(n10879), .A2(n5407), .ZN(n8430) );
  INV_X1 U5771 ( .A(n5409), .ZN(n5407) );
  INV_X1 U5772 ( .A(n7362), .ZN(n5417) );
  AND2_X1 U5773 ( .A1(n6414), .A2(n6402), .ZN(n6412) );
  AOI21_X1 U5774 ( .B1(n6373), .B2(n5262), .A(n5261), .ZN(n5260) );
  INV_X1 U5775 ( .A(n6051), .ZN(n5262) );
  INV_X1 U5776 ( .A(n6055), .ZN(n5261) );
  INV_X1 U5777 ( .A(n6373), .ZN(n5263) );
  INV_X1 U5778 ( .A(n5610), .ZN(n5609) );
  OAI21_X1 U5779 ( .B1(n5611), .B2(n6015), .A(n6014), .ZN(n5610) );
  NAND2_X1 U5780 ( .A1(n6255), .A2(n6011), .ZN(n5611) );
  NOR2_X1 U5781 ( .A1(n6015), .A2(n5613), .ZN(n5612) );
  INV_X1 U5782 ( .A(n6011), .ZN(n5613) );
  NAND2_X1 U5783 ( .A1(n6008), .A2(n9069), .ZN(n6011) );
  NAND2_X1 U5784 ( .A1(n9001), .A2(n6536), .ZN(n5683) );
  NOR2_X2 U5785 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5502) );
  INV_X1 U5786 ( .A(n5982), .ZN(n5586) );
  AND2_X1 U5787 ( .A1(n5978), .A2(n5976), .ZN(n5581) );
  NAND2_X1 U5788 ( .A1(n5622), .A2(n5625), .ZN(n5620) );
  AOI21_X1 U5789 ( .B1(n9279), .B2(n5167), .A(n5101), .ZN(n5239) );
  NAND2_X1 U5790 ( .A1(n8045), .A2(n5647), .ZN(n5646) );
  AND2_X1 U5791 ( .A1(n8827), .A2(n8828), .ZN(n5667) );
  AND2_X1 U5792 ( .A1(n6182), .A2(n7848), .ZN(n6199) );
  NAND2_X1 U5793 ( .A1(n5646), .A2(n5185), .ZN(n5642) );
  AND2_X1 U5794 ( .A1(n7959), .A2(n5648), .ZN(n5643) );
  INV_X1 U5795 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8669) );
  NAND2_X1 U5796 ( .A1(n9286), .A2(n5129), .ZN(n9345) );
  XNOR2_X1 U5797 ( .A(n7735), .B(n7930), .ZN(n7737) );
  AND2_X1 U5798 ( .A1(n5631), .A2(n9302), .ZN(n5627) );
  AOI21_X1 U5799 ( .B1(n5626), .B2(n5624), .A(n5623), .ZN(n5622) );
  INV_X1 U5800 ( .A(n5627), .ZN(n5624) );
  INV_X1 U5801 ( .A(n9358), .ZN(n5623) );
  INV_X1 U5802 ( .A(n5626), .ZN(n5625) );
  OR2_X1 U5803 ( .A1(n7306), .A2(n6524), .ZN(n7725) );
  OR2_X1 U5804 ( .A1(n6154), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6167) );
  AND2_X1 U5805 ( .A1(n5186), .A2(n8042), .ZN(n5369) );
  OR2_X1 U5806 ( .A1(n7352), .A2(n8355), .ZN(n7747) );
  OR2_X1 U5807 ( .A1(n5086), .A2(n7641), .ZN(n6104) );
  NAND4_X1 U5808 ( .A1(n6082), .A2(n6081), .A3(n6080), .A4(n6079), .ZN(n6098)
         );
  OR2_X1 U5809 ( .A1(n6470), .A2(n6078), .ZN(n6081) );
  OR2_X1 U5810 ( .A1(n5085), .A2(n7421), .ZN(n6088) );
  AND2_X1 U5811 ( .A1(n5473), .A2(n5472), .ZN(n7440) );
  NAND2_X1 U5812 ( .A1(n5871), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5472) );
  NOR2_X1 U5813 ( .A1(n5471), .A2(n10664), .ZN(n5470) );
  NOR2_X1 U5814 ( .A1(n7482), .A2(n5821), .ZN(n10680) );
  NOR2_X1 U5815 ( .A1(n10680), .A2(n10679), .ZN(n10678) );
  OR2_X1 U5816 ( .A1(n7479), .A2(n7480), .ZN(n5479) );
  AND3_X1 U5817 ( .A1(n5476), .A2(n5474), .A3(n5160), .ZN(n5875) );
  OR2_X1 U5818 ( .A1(n10715), .A2(n10716), .ZN(n5485) );
  AND3_X1 U5819 ( .A1(n5480), .A2(n5175), .A3(n5482), .ZN(n5880) );
  AND2_X1 U5820 ( .A1(n5924), .A2(n8130), .ZN(n8203) );
  NOR2_X1 U5821 ( .A1(n8499), .A2(n8500), .ZN(n8498) );
  NAND2_X1 U5822 ( .A1(n5491), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5490) );
  INV_X1 U5823 ( .A(n9417), .ZN(n5491) );
  NAND2_X1 U5824 ( .A1(n5229), .A2(n5226), .ZN(n5751) );
  AND4_X1 U5825 ( .A1(n5083), .A2(n5737), .A3(n5799), .A4(n5228), .ZN(n5226)
         );
  INV_X1 U5826 ( .A(n5798), .ZN(n5229) );
  INV_X1 U5827 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5228) );
  AND2_X1 U5828 ( .A1(n9424), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9426) );
  NAND2_X1 U5829 ( .A1(n5726), .A2(n5848), .ZN(n5566) );
  NOR2_X1 U5830 ( .A1(n9451), .A2(n5568), .ZN(n5567) );
  NOR2_X1 U5831 ( .A1(n9445), .A2(n9437), .ZN(n5494) );
  OAI21_X1 U5832 ( .B1(n9469), .B2(n5182), .A(n5572), .ZN(n9488) );
  INV_X1 U5833 ( .A(n9489), .ZN(n5573) );
  OR2_X1 U5834 ( .A1(n9469), .A2(n9468), .ZN(n5575) );
  INV_X1 U5835 ( .A(n5862), .ZN(n9512) );
  OR2_X1 U5836 ( .A1(n5859), .A2(n6297), .ZN(n5862) );
  AND2_X1 U5837 ( .A1(n9533), .A2(n6422), .ZN(n9281) );
  NAND2_X1 U5838 ( .A1(n5208), .A2(n5551), .ZN(n9574) );
  AOI21_X1 U5839 ( .B1(n5097), .B2(n5094), .A(n5143), .ZN(n5551) );
  NAND2_X1 U5840 ( .A1(n9599), .A2(n5097), .ZN(n5208) );
  NAND2_X1 U5841 ( .A1(n6362), .A2(n9349), .ZN(n6363) );
  AND2_X1 U5842 ( .A1(n6360), .A2(n6359), .ZN(n8820) );
  AOI21_X1 U5843 ( .B1(n9633), .B2(n9634), .A(n5192), .ZN(n9621) );
  NOR2_X1 U5844 ( .A1(n9719), .A2(n5193), .ZN(n5192) );
  NOR2_X1 U5845 ( .A1(n6338), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6349) );
  INV_X1 U5846 ( .A(n6287), .ZN(n6301) );
  NOR2_X1 U5847 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(n6301), .ZN(n6311) );
  NOR2_X1 U5848 ( .A1(n6288), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U5849 ( .A1(n8766), .A2(n6273), .ZN(n6288) );
  NAND2_X1 U5850 ( .A1(n8669), .A2(n6249), .ZN(n6261) );
  OR2_X1 U5851 ( .A1(n6212), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U5852 ( .A1(n8087), .A2(n6206), .ZN(n8094) );
  NAND2_X1 U5853 ( .A1(n7882), .A2(n7219), .ZN(n5500) );
  NAND2_X1 U5854 ( .A1(n5201), .A2(n6152), .ZN(n7919) );
  OR2_X1 U5855 ( .A1(n7760), .A2(n6151), .ZN(n5201) );
  INV_X1 U5856 ( .A(n5354), .ZN(n5353) );
  INV_X1 U5857 ( .A(n7680), .ZN(n5355) );
  NAND2_X1 U5858 ( .A1(n5199), .A2(n5197), .ZN(n7760) );
  AOI21_X1 U5859 ( .B1(n5200), .B2(n6126), .A(n5198), .ZN(n5197) );
  NAND2_X1 U5860 ( .A1(n7666), .A2(n5200), .ZN(n5199) );
  NOR2_X1 U5861 ( .A1(n9401), .A2(n7772), .ZN(n5198) );
  INV_X1 U5862 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9116) );
  NAND2_X1 U5863 ( .A1(n7680), .A2(n7200), .ZN(n7758) );
  NOR2_X1 U5864 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6141) );
  NAND2_X1 U5865 ( .A1(n5196), .A2(n6127), .ZN(n7683) );
  OR2_X1 U5866 ( .A1(n7666), .A2(n6126), .ZN(n5196) );
  CLKBUF_X1 U5867 ( .A(n7331), .Z(n7332) );
  AND2_X1 U5868 ( .A1(n6466), .A2(n8355), .ZN(n8292) );
  INV_X1 U5869 ( .A(n9635), .ZN(n9667) );
  INV_X1 U5870 ( .A(n9637), .ZN(n9668) );
  OR2_X1 U5871 ( .A1(n7306), .A2(n6523), .ZN(n8355) );
  NAND2_X1 U5872 ( .A1(n6405), .A2(n6404), .ZN(n8841) );
  NAND2_X1 U5873 ( .A1(n8122), .A2(n8262), .ZN(n8726) );
  AND2_X1 U5874 ( .A1(n5766), .A2(n5779), .ZN(n6488) );
  NAND2_X1 U5875 ( .A1(n5501), .A2(n5765), .ZN(n5762) );
  XNOR2_X1 U5876 ( .A(n5746), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7730) );
  NAND2_X1 U5877 ( .A1(n5745), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U5878 ( .A1(n5871), .A2(n5814), .ZN(n5816) );
  MUX2_X1 U5879 ( .A(n5815), .B(P2_IR_REG_31__SCAN_IN), .S(n5814), .Z(n5817)
         );
  NOR2_X1 U5880 ( .A1(n9813), .A2(n9812), .ZN(n9919) );
  AND2_X1 U5881 ( .A1(n9811), .A2(n9810), .ZN(n9812) );
  NAND2_X1 U5882 ( .A1(n9919), .A2(n9920), .ZN(n9918) );
  NOR2_X1 U5883 ( .A1(n6628), .A2(n10051), .ZN(n6627) );
  AOI21_X1 U5884 ( .B1(n5434), .B2(n9847), .A(n5135), .ZN(n5432) );
  AND2_X1 U5885 ( .A1(n5436), .A2(n5435), .ZN(n5434) );
  INV_X1 U5886 ( .A(n10026), .ZN(n5435) );
  OR2_X1 U5887 ( .A1(n9847), .A2(n9848), .ZN(n5436) );
  INV_X1 U5888 ( .A(n9823), .ZN(n9998) );
  AND2_X1 U5889 ( .A1(n9882), .A2(n9880), .ZN(n10015) );
  NAND2_X1 U5890 ( .A1(n7516), .A2(n5272), .ZN(n7518) );
  NAND2_X1 U5891 ( .A1(n9953), .A2(n7973), .ZN(n5272) );
  INV_X1 U5892 ( .A(n9860), .ZN(n7647) );
  NAND2_X1 U5893 ( .A1(n5428), .A2(n5132), .ZN(n10048) );
  AND2_X1 U5894 ( .A1(n9838), .A2(n9837), .ZN(n9843) );
  INV_X1 U5895 ( .A(n8070), .ZN(n8068) );
  MUX2_X1 U5896 ( .A(n6976), .B(n6975), .S(n7033), .Z(n6983) );
  AND4_X1 U5897 ( .A1(n6798), .A2(n6797), .A3(n6796), .A4(n6795), .ZN(n8746)
         );
  AND4_X1 U5898 ( .A1(n6779), .A2(n6778), .A3(n6777), .A4(n6776), .ZN(n8372)
         );
  NOR2_X1 U5899 ( .A1(n7589), .A2(n5114), .ZN(n10766) );
  NOR2_X1 U5900 ( .A1(n10766), .A2(n10765), .ZN(n10764) );
  NAND2_X1 U5901 ( .A1(n7874), .A2(n7875), .ZN(n8215) );
  OR2_X1 U5902 ( .A1(n8591), .A2(n8590), .ZN(n5421) );
  AND2_X1 U5903 ( .A1(n10140), .A2(n10158), .ZN(n10169) );
  AND2_X1 U5904 ( .A1(n10181), .A2(n5418), .ZN(n10183) );
  NAND2_X1 U5905 ( .A1(n10182), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5418) );
  NAND2_X1 U5906 ( .A1(n10487), .A2(n5411), .ZN(n5410) );
  INV_X1 U5907 ( .A(n5412), .ZN(n5411) );
  OR2_X1 U5908 ( .A1(n10320), .A2(n5413), .ZN(n10285) );
  NAND2_X1 U5909 ( .A1(n10298), .A2(n5190), .ZN(n10284) );
  OR2_X1 U5910 ( .A1(n10270), .A2(n10501), .ZN(n5190) );
  INV_X1 U5911 ( .A(n10351), .ZN(n10318) );
  NAND2_X1 U5912 ( .A1(n10362), .A2(n10239), .ZN(n5512) );
  AND2_X1 U5913 ( .A1(n10241), .A2(n5514), .ZN(n5513) );
  AND2_X1 U5914 ( .A1(n10393), .A2(n5150), .ZN(n10330) );
  AND2_X1 U5915 ( .A1(n6997), .A2(n10242), .ZN(n10334) );
  NAND2_X1 U5916 ( .A1(n10393), .A2(n5391), .ZN(n10343) );
  NAND2_X1 U5917 ( .A1(n10377), .A2(n10238), .ZN(n10361) );
  NAND2_X1 U5918 ( .A1(n10361), .A2(n10362), .ZN(n10360) );
  NAND2_X1 U5919 ( .A1(n10368), .A2(n5118), .ZN(n10356) );
  NAND2_X1 U5920 ( .A1(n10393), .A2(n10376), .ZN(n10371) );
  NAND2_X1 U5921 ( .A1(n10370), .A2(n10369), .ZN(n10368) );
  OR2_X1 U5922 ( .A1(n6882), .A2(n6881), .ZN(n6900) );
  INV_X1 U5923 ( .A(n5688), .ZN(n5687) );
  OAI21_X1 U5924 ( .B1(n5690), .B2(n7017), .A(n5716), .ZN(n5688) );
  AND4_X1 U5925 ( .A1(n6887), .A2(n6886), .A3(n6885), .A4(n6884), .ZN(n10463)
         );
  NAND2_X1 U5926 ( .A1(n8644), .A2(n10975), .ZN(n10555) );
  NAND2_X1 U5927 ( .A1(n8550), .A2(n7015), .ZN(n8639) );
  NAND2_X1 U5928 ( .A1(n6827), .A2(n6826), .ZN(n9799) );
  INV_X1 U5929 ( .A(n5525), .ZN(n5524) );
  OAI21_X1 U5930 ( .B1(n5527), .B2(n5526), .A(n10940), .ZN(n5525) );
  AOI21_X1 U5931 ( .B1(n8555), .B2(n5674), .A(n5138), .ZN(n5673) );
  INV_X1 U5932 ( .A(n8428), .ZN(n5674) );
  NOR2_X1 U5933 ( .A1(n6775), .A2(n6763), .ZN(n6791) );
  NOR2_X1 U5934 ( .A1(n10879), .A2(n8345), .ZN(n8378) );
  AOI21_X1 U5935 ( .B1(n10890), .B2(n5679), .A(n5141), .ZN(n5678) );
  INV_X1 U5936 ( .A(n8274), .ZN(n5679) );
  OR2_X1 U5937 ( .A1(n10878), .A2(n10899), .ZN(n10879) );
  INV_X1 U5938 ( .A(n5535), .ZN(n5534) );
  INV_X1 U5939 ( .A(n5532), .ZN(n5533) );
  AOI21_X1 U5940 ( .B1(n7088), .B2(n7003), .A(n5536), .ZN(n5535) );
  AND2_X1 U5941 ( .A1(n8022), .A2(n8002), .ZN(n8189) );
  NOR2_X1 U5942 ( .A1(n10814), .A2(n8072), .ZN(n8022) );
  OR2_X1 U5943 ( .A1(n10813), .A2(n10829), .ZN(n10814) );
  NAND2_X1 U5944 ( .A1(n10785), .A2(n7806), .ZN(n10813) );
  NOR2_X1 U5945 ( .A1(n10784), .A2(n10795), .ZN(n10785) );
  NOR2_X1 U5946 ( .A1(n7973), .A2(n7977), .ZN(n7970) );
  INV_X1 U5947 ( .A(n11022), .ZN(n11027) );
  NAND2_X1 U5948 ( .A1(n8426), .A2(n8425), .ZN(n5675) );
  INV_X1 U5949 ( .A(n10557), .ZN(n11031) );
  OAI21_X1 U5950 ( .B1(n10574), .B2(P1_D_REG_0__SCAN_IN), .A(n10576), .ZN(
        n7946) );
  AND2_X1 U5951 ( .A1(n7948), .A2(n7538), .ZN(n7552) );
  INV_X1 U5952 ( .A(n7976), .ZN(n7977) );
  XNOR2_X1 U5953 ( .A(n6548), .B(n6547), .ZN(n6549) );
  NAND2_X1 U5954 ( .A1(n5700), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6556) );
  AND2_X1 U5955 ( .A1(n5705), .A2(n5702), .ZN(n5701) );
  XNOR2_X1 U5956 ( .A(n6413), .B(n6412), .ZN(n8755) );
  AND2_X1 U5957 ( .A1(n6553), .A2(n5704), .ZN(n5703) );
  INV_X1 U5958 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5704) );
  XNOR2_X1 U5959 ( .A(n6384), .B(n6383), .ZN(n8632) );
  NAND2_X1 U5960 ( .A1(n5259), .A2(n5260), .ZN(n6384) );
  OR2_X1 U5961 ( .A1(n6067), .A2(n5263), .ZN(n5259) );
  XNOR2_X1 U5962 ( .A(n7159), .B(P1_IR_REG_24__SCAN_IN), .ZN(n7492) );
  NAND2_X1 U5963 ( .A1(n6545), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6546) );
  INV_X1 U5964 ( .A(n5589), .ZN(n5588) );
  OAI21_X1 U5965 ( .B1(n5592), .B2(n5590), .A(n6035), .ZN(n5589) );
  NAND2_X1 U5966 ( .A1(n5591), .A2(n6029), .ZN(n5590) );
  AND2_X1 U5967 ( .A1(n6039), .A2(n6038), .ZN(n6332) );
  NAND2_X1 U5968 ( .A1(n6893), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6540) );
  NAND2_X1 U5969 ( .A1(n6026), .A2(n6025), .ZN(n6308) );
  NAND2_X1 U5970 ( .A1(n6542), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6850) );
  NAND2_X1 U5971 ( .A1(n5250), .A2(n5615), .ZN(n6232) );
  OAI21_X1 U5972 ( .B1(n6207), .B2(n5995), .A(n5997), .ZN(n6221) );
  AND2_X1 U5973 ( .A1(n6741), .A2(n6808), .ZN(n7873) );
  AND2_X1 U5974 ( .A1(n6716), .A2(n6715), .ZN(n7620) );
  XNOR2_X1 U5975 ( .A(n5979), .B(n9083), .ZN(n6148) );
  NAND2_X1 U5976 ( .A1(n5977), .A2(n5976), .ZN(n6136) );
  CLKBUF_X1 U5977 ( .A(n6689), .Z(n6690) );
  XNOR2_X1 U5978 ( .A(n5968), .B(SI_1_), .ZN(n6084) );
  NOR2_X1 U5979 ( .A1(n7297), .A2(n5302), .ZN(n5301) );
  INV_X1 U5980 ( .A(n9579), .ZN(n5302) );
  NAND2_X1 U5981 ( .A1(n5644), .A2(n5643), .ZN(n8046) );
  NOR2_X1 U5982 ( .A1(n5652), .A2(n9355), .ZN(n5650) );
  NOR2_X1 U5983 ( .A1(n5653), .A2(n5656), .ZN(n5652) );
  NOR2_X1 U5984 ( .A1(n5659), .A2(n5167), .ZN(n5656) );
  NAND2_X1 U5985 ( .A1(n5654), .A2(n5658), .ZN(n5651) );
  NAND2_X1 U5986 ( .A1(n5655), .A2(n9279), .ZN(n5654) );
  NAND2_X1 U5987 ( .A1(n5218), .A2(n5632), .ZN(n8709) );
  NAND2_X1 U5988 ( .A1(n5217), .A2(n5635), .ZN(n5218) );
  NAND2_X1 U5989 ( .A1(n5666), .A2(n7742), .ZN(n7765) );
  NAND2_X1 U5990 ( .A1(n9271), .A2(n9270), .ZN(n9269) );
  NAND2_X1 U5991 ( .A1(n8046), .A2(n5646), .ZN(n8110) );
  NAND2_X1 U5992 ( .A1(n7936), .A2(n7935), .ZN(n7934) );
  AND4_X1 U5993 ( .A1(n6343), .A2(n6342), .A3(n6341), .A4(n6340), .ZN(n9636)
         );
  NAND2_X1 U5994 ( .A1(n9288), .A2(n9287), .ZN(n9286) );
  NAND2_X1 U5995 ( .A1(n5663), .A2(n5661), .ZN(n8057) );
  NAND2_X1 U5996 ( .A1(n5662), .A2(n7777), .ZN(n5661) );
  NAND2_X1 U5997 ( .A1(n9306), .A2(n9302), .ZN(n5630) );
  INV_X1 U5998 ( .A(n9295), .ZN(n9325) );
  NAND2_X1 U5999 ( .A1(n7777), .A2(n5209), .ZN(n7767) );
  NAND2_X1 U6000 ( .A1(n5210), .A2(n9401), .ZN(n5209) );
  AND2_X1 U6001 ( .A1(n7765), .A2(n5660), .ZN(n7778) );
  INV_X1 U6002 ( .A(n5662), .ZN(n5660) );
  NAND2_X1 U6003 ( .A1(n7765), .A2(n5665), .ZN(n7768) );
  NAND2_X1 U6004 ( .A1(n5639), .A2(n5213), .ZN(n8113) );
  INV_X1 U6005 ( .A(n5640), .ZN(n5639) );
  NAND2_X1 U6006 ( .A1(n7956), .A2(n5641), .ZN(n5213) );
  OAI21_X1 U6007 ( .B1(n5643), .B2(n5642), .A(n8109), .ZN(n5640) );
  NAND2_X1 U6008 ( .A1(n7750), .A2(n7749), .ZN(n9328) );
  NAND2_X1 U6009 ( .A1(n5636), .A2(n5635), .ZN(n8708) );
  AND2_X1 U6010 ( .A1(n5636), .A2(n5117), .ZN(n8665) );
  NAND2_X1 U6011 ( .A1(n8664), .A2(n8663), .ZN(n5636) );
  NAND2_X1 U6012 ( .A1(n9286), .A2(n8819), .ZN(n9347) );
  NAND2_X1 U6013 ( .A1(n5225), .A2(n5712), .ZN(n8470) );
  OR2_X1 U6014 ( .A1(n8437), .A2(n9396), .ZN(n5225) );
  INV_X1 U6015 ( .A(n5621), .ZN(n9359) );
  AOI21_X1 U6016 ( .B1(n9306), .B2(n5627), .A(n5625), .ZN(n5621) );
  OAI21_X1 U6017 ( .B1(n9306), .B2(n5625), .A(n5622), .ZN(n9357) );
  INV_X1 U6018 ( .A(n5214), .ZN(n8055) );
  AND2_X1 U6019 ( .A1(n8764), .A2(n8761), .ZN(n8762) );
  XNOR2_X1 U6020 ( .A(n5752), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7354) );
  OR2_X1 U6021 ( .A1(n5501), .A2(n5806), .ZN(n5752) );
  INV_X1 U6022 ( .A(n5278), .ZN(n5275) );
  NOR2_X1 U6023 ( .A1(n5095), .A2(n8042), .ZN(n5274) );
  AOI21_X1 U6024 ( .B1(n5278), .B2(n8042), .A(n5277), .ZN(n5276) );
  NAND2_X1 U6025 ( .A1(n5370), .A2(n5375), .ZN(n5277) );
  INV_X1 U6026 ( .A(n8415), .ZN(n5375) );
  NAND2_X1 U6027 ( .A1(n7329), .A2(n5120), .ZN(n5370) );
  OR2_X1 U6028 ( .A1(n5599), .A2(n6480), .ZN(n5371) );
  INV_X1 U6029 ( .A(n9589), .ZN(n9386) );
  INV_X1 U6030 ( .A(n9638), .ZN(n9611) );
  AND4_X1 U6031 ( .A1(n6204), .A2(n6203), .A3(n6202), .A4(n6201), .ZN(n8449)
         );
  CLKBUF_X1 U6032 ( .A(n6098), .Z(n9404) );
  OR2_X1 U6033 ( .A1(n7722), .A2(n5942), .ZN(n10657) );
  NAND2_X1 U6034 ( .A1(n5870), .A2(n5869), .ZN(n10665) );
  NAND2_X1 U6035 ( .A1(n5474), .A2(n5476), .ZN(n10675) );
  NOR2_X1 U6036 ( .A1(n10696), .A2(n5824), .ZN(n7463) );
  NOR2_X1 U6037 ( .A1(n8200), .A2(n8199), .ZN(n8198) );
  NOR2_X1 U6038 ( .A1(n8126), .A2(n5838), .ZN(n8208) );
  NOR2_X1 U6039 ( .A1(n8496), .A2(n8497), .ZN(n8495) );
  NAND2_X1 U6040 ( .A1(n5176), .A2(n5496), .ZN(n5495) );
  OR2_X1 U6041 ( .A1(n9460), .A2(n5891), .ZN(n5460) );
  INV_X1 U6042 ( .A(n5388), .ZN(n5379) );
  OAI21_X1 U6043 ( .B1(n9553), .B2(n9653), .A(n9552), .ZN(n9687) );
  OAI22_X1 U6044 ( .A1(n9576), .A2(n9635), .B1(n9637), .B2(n9550), .ZN(n9551)
         );
  NAND2_X1 U6045 ( .A1(n9565), .A2(n9564), .ZN(n9690) );
  INV_X1 U6046 ( .A(n9563), .ZN(n9564) );
  NAND2_X1 U6047 ( .A1(n9562), .A2(n9664), .ZN(n9565) );
  NAND2_X1 U6048 ( .A1(n9696), .A2(n6462), .ZN(n9567) );
  AND2_X1 U6049 ( .A1(n5960), .A2(n6419), .ZN(n9577) );
  OR2_X1 U6050 ( .A1(n9599), .A2(n5094), .ZN(n5552) );
  NAND2_X1 U6051 ( .A1(n5359), .A2(n7167), .ZN(n9603) );
  NAND2_X1 U6052 ( .A1(n9626), .A2(n7168), .ZN(n9615) );
  INV_X1 U6053 ( .A(n8820), .ZN(n9714) );
  OR2_X1 U6054 ( .A1(n6460), .A2(n5468), .ZN(n5464) );
  NAND2_X1 U6055 ( .A1(n9663), .A2(n6331), .ZN(n9651) );
  NAND2_X1 U6056 ( .A1(n6337), .A2(n6336), .ZN(n9657) );
  NAND2_X1 U6057 ( .A1(n6323), .A2(n6322), .ZN(n9674) );
  NAND2_X1 U6058 ( .A1(n5548), .A2(n5549), .ZN(n8695) );
  OR2_X1 U6059 ( .A1(n6294), .A2(n6458), .ZN(n5548) );
  NAND2_X1 U6060 ( .A1(n8722), .A2(n6459), .ZN(n8700) );
  NAND2_X1 U6061 ( .A1(n6299), .A2(n6298), .ZN(n9321) );
  NAND2_X1 U6062 ( .A1(n6285), .A2(n6284), .ZN(n9312) );
  NAND2_X1 U6063 ( .A1(n6271), .A2(n6270), .ZN(n8760) );
  NAND2_X1 U6064 ( .A1(n5537), .A2(n5542), .ZN(n8627) );
  NAND2_X1 U6065 ( .A1(n8458), .A2(n6266), .ZN(n5537) );
  NAND2_X1 U6066 ( .A1(n8456), .A2(n6266), .ZN(n8533) );
  NAND2_X1 U6067 ( .A1(n6259), .A2(n6258), .ZN(n8706) );
  OAI21_X1 U6068 ( .B1(n8268), .B2(n8266), .A(n7240), .ZN(n8462) );
  INV_X1 U6069 ( .A(n8471), .ZN(n8524) );
  NAND2_X1 U6070 ( .A1(n8088), .A2(n5205), .ZN(n5202) );
  NAND2_X1 U6071 ( .A1(n8096), .A2(n6219), .ZN(n8323) );
  NAND2_X1 U6072 ( .A1(n7665), .A2(n7667), .ZN(n7664) );
  NAND2_X1 U6073 ( .A1(n6450), .A2(n7191), .ZN(n7665) );
  INV_X1 U6074 ( .A(n9677), .ZN(n9629) );
  OR2_X1 U6075 ( .A1(n8358), .A2(n9592), .ZN(n9647) );
  INV_X1 U6076 ( .A(n9647), .ZN(n10869) );
  OR2_X1 U6077 ( .A1(n7301), .A2(n7368), .ZN(n6124) );
  INV_X2 U6078 ( .A(n9735), .ZN(n9683) );
  INV_X1 U6079 ( .A(n7328), .ZN(n9741) );
  AOI21_X1 U6080 ( .B1(n9258), .B2(n7308), .A(n7302), .ZN(n9744) );
  NOR2_X1 U6081 ( .A1(n9687), .A2(n9686), .ZN(n9745) );
  AND2_X1 U6082 ( .A1(n9685), .A2(n9733), .ZN(n9686) );
  INV_X1 U6083 ( .A(n8841), .ZN(n9752) );
  AND2_X1 U6084 ( .A1(n6063), .A2(n6062), .ZN(n9756) );
  INV_X1 U6085 ( .A(n6393), .ZN(n9760) );
  AND2_X1 U6086 ( .A1(n6376), .A2(n6375), .ZN(n9764) );
  AND2_X1 U6087 ( .A1(n6180), .A2(n6179), .ZN(n8514) );
  AND2_X1 U6088 ( .A1(n6176), .A2(n6175), .ZN(n7968) );
  INV_X1 U6089 ( .A(n11017), .ZN(n11015) );
  AND2_X1 U6090 ( .A1(n7721), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8783) );
  INV_X1 U6091 ( .A(n6488), .ZN(n8784) );
  XNOR2_X1 U6092 ( .A(n5757), .B(n5756), .ZN(n6485) );
  NAND2_X1 U6093 ( .A1(n5755), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5757) );
  XNOR2_X1 U6094 ( .A(n5759), .B(n5758), .ZN(n6484) );
  INV_X1 U6095 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8264) );
  INV_X1 U6096 ( .A(n7354), .ZN(n8262) );
  INV_X1 U6097 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8044) );
  INV_X1 U6098 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7819) );
  INV_X1 U6099 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7700) );
  INV_X1 U6100 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7557) );
  NOR2_X1 U6101 ( .A1(n5798), .A2(n5230), .ZN(n5796) );
  NAND2_X1 U6102 ( .A1(n5083), .A2(n5799), .ZN(n5230) );
  INV_X1 U6103 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7399) );
  INV_X1 U6104 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7393) );
  INV_X1 U6105 ( .A(n10686), .ZN(n7369) );
  NAND2_X1 U6106 ( .A1(n5817), .A2(n5816), .ZN(n7363) );
  NAND2_X1 U6107 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5457) );
  NAND2_X1 U6108 ( .A1(n6600), .A2(n6599), .ZN(n10520) );
  INV_X1 U6109 ( .A(n9892), .ZN(n5282) );
  AND2_X1 U6110 ( .A1(n9911), .A2(n5280), .ZN(n5279) );
  NAND2_X1 U6111 ( .A1(n9892), .A2(n5281), .ZN(n5280) );
  AND2_X1 U6112 ( .A1(n9904), .A2(n9903), .ZN(n9966) );
  NAND2_X1 U6113 ( .A1(n6586), .A2(n6585), .ZN(n10495) );
  NAND2_X1 U6114 ( .A1(n5433), .A2(n5432), .ZN(n9975) );
  NAND2_X1 U6115 ( .A1(n9937), .A2(n5434), .ZN(n5433) );
  NAND2_X1 U6116 ( .A1(n6609), .A2(n6608), .ZN(n10531) );
  NAND2_X1 U6117 ( .A1(n5254), .A2(n8740), .ZN(n8744) );
  NAND2_X1 U6118 ( .A1(n5447), .A2(n7829), .ZN(n7838) );
  NAND2_X1 U6119 ( .A1(n8329), .A2(n8328), .ZN(n5439) );
  AOI21_X1 U6120 ( .B1(n9937), .B2(n9848), .A(n9847), .ZN(n10025) );
  NAND2_X1 U6121 ( .A1(n9803), .A2(n9802), .ZN(n10036) );
  AND4_X1 U6122 ( .A1(n6614), .A2(n6613), .A3(n6612), .A4(n6611), .ZN(n10263)
         );
  NAND2_X1 U6123 ( .A1(n8795), .A2(n8796), .ZN(n8794) );
  INV_X1 U6124 ( .A(n9843), .ZN(n10058) );
  AND2_X1 U6125 ( .A1(n5449), .A2(n8147), .ZN(n8159) );
  NAND2_X1 U6126 ( .A1(n6940), .A2(n6939), .ZN(n10506) );
  AND2_X1 U6127 ( .A1(n7811), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10071) );
  NOR2_X1 U6128 ( .A1(n10041), .A2(n10462), .ZN(n10087) );
  AND2_X1 U6129 ( .A1(n7524), .A2(n7523), .ZN(n10081) );
  AND4_X1 U6130 ( .A1(n6817), .A2(n6816), .A3(n6815), .A4(n6814), .ZN(n10094)
         );
  OR2_X1 U6131 ( .A1(n7511), .A2(n7359), .ZN(n10104) );
  INV_X1 U6132 ( .A(n7562), .ZN(n10654) );
  NOR2_X1 U6133 ( .A1(n10764), .A2(n5424), .ZN(n7604) );
  NOR2_X1 U6134 ( .A1(n7572), .A2(n5425), .ZN(n5424) );
  NOR2_X1 U6135 ( .A1(n7604), .A2(n7603), .ZN(n7602) );
  NOR2_X1 U6136 ( .A1(n7701), .A2(n5169), .ZN(n7704) );
  NOR2_X1 U6137 ( .A1(n7704), .A2(n7703), .ZN(n7872) );
  OR2_X1 U6138 ( .A1(n8216), .A2(n5423), .ZN(n10110) );
  INV_X1 U6139 ( .A(n10112), .ZN(n5423) );
  INV_X1 U6140 ( .A(n8216), .ZN(n10111) );
  AND2_X1 U6141 ( .A1(n10110), .A2(n5422), .ZN(n8219) );
  NAND2_X1 U6142 ( .A1(n10105), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5422) );
  INV_X1 U6143 ( .A(n5421), .ZN(n10123) );
  NAND2_X1 U6144 ( .A1(n5421), .A2(n5420), .ZN(n10125) );
  NAND2_X1 U6145 ( .A1(n10124), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6146 ( .A1(n10125), .A2(n10126), .ZN(n10138) );
  INV_X1 U6147 ( .A(n10222), .ZN(n10763) );
  INV_X1 U6148 ( .A(n10226), .ZN(n10487) );
  AOI21_X1 U6149 ( .B1(n10271), .B2(n10550), .A(n10251), .ZN(n10252) );
  XNOR2_X1 U6150 ( .A(n5523), .B(n10248), .ZN(n10253) );
  NOR2_X1 U6151 ( .A1(n10301), .A2(n10246), .ZN(n10292) );
  INV_X1 U6152 ( .A(n10495), .ZN(n10290) );
  AND2_X1 U6153 ( .A1(n6955), .A2(n6954), .ZN(n10308) );
  NAND2_X1 U6154 ( .A1(n10313), .A2(n5722), .ZN(n10300) );
  INV_X1 U6155 ( .A(n10506), .ZN(n10326) );
  INV_X1 U6156 ( .A(n10520), .ZN(n10265) );
  NAND2_X1 U6157 ( .A1(n5696), .A2(n5695), .ZN(n10529) );
  AND2_X1 U6158 ( .A1(n10391), .A2(n5096), .ZN(n5695) );
  AND2_X1 U6159 ( .A1(n5694), .A2(n5096), .ZN(n10392) );
  INV_X1 U6160 ( .A(n5694), .ZN(n10400) );
  NAND2_X1 U6161 ( .A1(n6635), .A2(n6634), .ZN(n10428) );
  AND2_X1 U6162 ( .A1(n10461), .A2(n7104), .ZN(n10448) );
  OR2_X1 U6163 ( .A1(n10546), .A2(n5690), .ZN(n10468) );
  NOR2_X1 U6164 ( .A1(n10546), .A2(n5692), .ZN(n10470) );
  NAND2_X1 U6165 ( .A1(n5508), .A2(n5509), .ZN(n10549) );
  OR2_X1 U6166 ( .A1(n11005), .A2(n7952), .ZN(n10995) );
  NAND2_X1 U6167 ( .A1(n7009), .A2(n7008), .ZN(n8421) );
  NAND2_X1 U6168 ( .A1(n10573), .A2(n7526), .ZN(n10472) );
  NAND2_X1 U6169 ( .A1(n8273), .A2(n8272), .ZN(n5681) );
  INV_X1 U6170 ( .A(n10995), .ZN(n10956) );
  INV_X1 U6171 ( .A(n10472), .ZN(n10992) );
  AND2_X2 U6172 ( .A1(n7552), .A2(n7539), .ZN(n11037) );
  NAND2_X1 U6173 ( .A1(n5267), .A2(n5264), .ZN(n5271) );
  NAND2_X1 U6174 ( .A1(n6560), .A2(n5516), .ZN(n10580) );
  NOR2_X1 U6175 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n5516) );
  NAND2_X1 U6176 ( .A1(n5404), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6555) );
  INV_X1 U6177 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9148) );
  INV_X1 U6178 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n9154) );
  INV_X1 U6179 ( .A(n7492), .ZN(n8587) );
  INV_X1 U6180 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9156) );
  INV_X1 U6181 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8084) );
  INV_X1 U6182 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8041) );
  CLKBUF_X1 U6183 ( .A(n7507), .Z(n10219) );
  NAND2_X1 U6184 ( .A1(n6867), .A2(n6538), .ZN(n6891) );
  INV_X1 U6185 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7559) );
  INV_X1 U6186 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9180) );
  INV_X1 U6187 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7396) );
  INV_X1 U6188 ( .A(n6704), .ZN(n7388) );
  XNOR2_X1 U6189 ( .A(n5426), .B(P1_IR_REG_1__SCAN_IN), .ZN(n7562) );
  NOR2_X1 U6190 ( .A1(n6838), .A2(n5427), .ZN(n5426) );
  INV_X1 U6191 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10736) );
  AOI21_X1 U6192 ( .B1(n7294), .B2(n5301), .A(n5299), .ZN(n5295) );
  NAND2_X1 U6193 ( .A1(n5234), .A2(n5658), .ZN(n5233) );
  NOR2_X1 U6194 ( .A1(n10712), .A2(n5829), .ZN(n7847) );
  OR2_X1 U6195 ( .A1(n9504), .A2(n5576), .ZN(P2_U3199) );
  OAI211_X1 U6196 ( .C1(n9508), .C2(n10717), .A(n5578), .B(n5577), .ZN(n5576)
         );
  NOR2_X1 U6197 ( .A1(n9511), .A2(n5140), .ZN(n9503) );
  AND2_X1 U6198 ( .A1(n9530), .A2(n9529), .ZN(n9531) );
  OR2_X1 U6199 ( .A1(n5950), .A2(n5949), .ZN(P2_U3201) );
  NAND2_X1 U6200 ( .A1(n6517), .A2(n9735), .ZN(n6532) );
  OAI21_X1 U6201 ( .B1(n7149), .B2(n7508), .A(n7148), .ZN(n7165) );
  INV_X1 U6202 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7909) );
  AND2_X1 U6203 ( .A1(n5554), .A2(n6331), .ZN(n5093) );
  AND2_X1 U6204 ( .A1(n9764), .A2(n9588), .ZN(n5094) );
  AND2_X1 U6205 ( .A1(n7329), .A2(n5105), .ZN(n5095) );
  OR2_X1 U6206 ( .A1(n10537), .A2(n5699), .ZN(n5096) );
  INV_X1 U6207 ( .A(n5249), .ZN(n5248) );
  NAND2_X1 U6208 ( .A1(n5615), .A2(n6231), .ZN(n5249) );
  INV_X1 U6209 ( .A(n9601), .ZN(n9622) );
  AND4_X1 U6210 ( .A1(n6077), .A2(n6076), .A3(n6075), .A4(n6074), .ZN(n9601)
         );
  INV_X1 U6211 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5954) );
  AND2_X1 U6212 ( .A1(n5112), .A2(n6394), .ZN(n5097) );
  AND2_X1 U6213 ( .A1(n5458), .A2(n5187), .ZN(n5098) );
  INV_X1 U6214 ( .A(n7986), .ZN(n5536) );
  AND2_X1 U6215 ( .A1(n7267), .A2(n5465), .ZN(n5099) );
  OR3_X1 U6216 ( .A1(n7139), .A2(n7161), .A3(n7525), .ZN(n5100) );
  AND2_X1 U6217 ( .A1(n9278), .A2(n9385), .ZN(n5101) );
  AND2_X1 U6218 ( .A1(n5236), .A2(n5116), .ZN(n5102) );
  INV_X1 U6219 ( .A(n9676), .ZN(n6330) );
  AND2_X1 U6220 ( .A1(n7265), .A2(n7258), .ZN(n9676) );
  INV_X1 U6221 ( .A(n5111), .ZN(n5614) );
  INV_X1 U6222 ( .A(n10537), .ZN(n10407) );
  NAND2_X1 U6223 ( .A1(n6616), .A2(n6615), .ZN(n10537) );
  NAND2_X1 U6224 ( .A1(n6347), .A2(n6346), .ZN(n9719) );
  AND2_X1 U6225 ( .A1(n5609), .A2(n5607), .ZN(n5103) );
  INV_X1 U6226 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5806) );
  INV_X1 U6227 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9236) );
  INV_X1 U6228 ( .A(n6689), .ZN(n5283) );
  NAND2_X1 U6229 ( .A1(n8468), .A2(n8473), .ZN(n5104) );
  AND2_X1 U6230 ( .A1(n7330), .A2(n5186), .ZN(n5105) );
  AND2_X1 U6231 ( .A1(n5775), .A2(n5562), .ZN(n5106) );
  AND2_X1 U6232 ( .A1(n5260), .A2(n6383), .ZN(n5107) );
  NAND2_X1 U6233 ( .A1(n5543), .A2(n7340), .ZN(n8456) );
  OR2_X1 U6234 ( .A1(n6535), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5108) );
  INV_X1 U6235 ( .A(n9355), .ZN(n5658) );
  INV_X1 U6236 ( .A(n5191), .ZN(n7353) );
  NAND4_X1 U6237 ( .A1(n6653), .A2(n6652), .A3(n6651), .A4(n6650), .ZN(n7973)
         );
  INV_X1 U6238 ( .A(n6692), .ZN(n6895) );
  NAND2_X2 U6239 ( .A1(n5959), .A2(n5958), .ZN(n6102) );
  INV_X1 U6240 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6838) );
  NAND2_X1 U6241 ( .A1(n6988), .A2(n5403), .ZN(n7152) );
  INV_X1 U6242 ( .A(n10099), .ZN(n5344) );
  OR2_X1 U6243 ( .A1(n10320), .A2(n5410), .ZN(n5109) );
  INV_X1 U6244 ( .A(n5452), .ZN(n7509) );
  NAND2_X1 U6245 ( .A1(n7146), .A2(n5287), .ZN(n5452) );
  INV_X1 U6246 ( .A(n8149), .ZN(n8002) );
  AND2_X1 U6247 ( .A1(n9918), .A2(n9814), .ZN(n5110) );
  INV_X1 U6248 ( .A(n7467), .ZN(n7374) );
  XNOR2_X1 U6249 ( .A(n5825), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7467) );
  OR2_X1 U6250 ( .A1(n6220), .A2(n5617), .ZN(n5111) );
  NAND2_X1 U6251 ( .A1(n9334), .A2(n9612), .ZN(n5112) );
  AND2_X1 U6252 ( .A1(n5740), .A2(n5216), .ZN(n5113) );
  OR2_X1 U6253 ( .A1(n10543), .A2(n10463), .ZN(n7107) );
  INV_X1 U6254 ( .A(n9618), .ZN(n9710) );
  AND2_X1 U6255 ( .A1(n6070), .A2(n6069), .ZN(n9618) );
  NAND2_X1 U6256 ( .A1(n10102), .A2(n10816), .ZN(n7046) );
  AND2_X1 U6257 ( .A1(n7595), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5114) );
  INV_X1 U6258 ( .A(n8555), .ZN(n5528) );
  XNOR2_X1 U6259 ( .A(n5271), .B(n6981), .ZN(n7309) );
  NAND2_X1 U6260 ( .A1(n5211), .A2(n8058), .ZN(n7777) );
  INV_X1 U6261 ( .A(n6174), .ZN(n5984) );
  XNOR2_X1 U6262 ( .A(n5985), .B(SI_7_), .ZN(n6174) );
  XOR2_X1 U6263 ( .A(n6084), .B(n6083), .Z(n5115) );
  OR2_X1 U6264 ( .A1(n9280), .A2(n5235), .ZN(n5116) );
  AND2_X1 U6265 ( .A1(n7218), .A2(n7225), .ZN(n8086) );
  XNOR2_X1 U6266 ( .A(n9555), .B(n10659), .ZN(n9548) );
  INV_X1 U6267 ( .A(n9548), .ZN(n9556) );
  INV_X1 U6268 ( .A(n7258), .ZN(n5466) );
  NAND2_X1 U6269 ( .A1(n6925), .A2(n6924), .ZN(n10510) );
  INV_X1 U6270 ( .A(n10510), .ZN(n5390) );
  NAND2_X1 U6271 ( .A1(n9262), .A2(n8827), .ZN(n9324) );
  NAND2_X1 U6272 ( .A1(n8662), .A2(n9394), .ZN(n5117) );
  INV_X1 U6273 ( .A(n9602), .ZN(n9387) );
  AND4_X1 U6274 ( .A1(n6392), .A2(n6391), .A3(n6390), .A4(n6389), .ZN(n9602)
         );
  INV_X1 U6275 ( .A(n5488), .ZN(n7667) );
  NAND2_X1 U6276 ( .A1(n7213), .A2(n7199), .ZN(n5488) );
  INV_X1 U6277 ( .A(n8186), .ZN(n8272) );
  XNOR2_X1 U6278 ( .A(n10858), .B(n5344), .ZN(n8186) );
  NAND2_X1 U6279 ( .A1(n6992), .A2(n10245), .ZN(n10302) );
  INV_X1 U6280 ( .A(n10302), .ZN(n5522) );
  OR2_X1 U6281 ( .A1(n10376), .A2(n10264), .ZN(n5118) );
  OR2_X1 U6282 ( .A1(n7734), .A2(n9404), .ZN(n5119) );
  AND2_X1 U6283 ( .A1(n7330), .A2(n5369), .ZN(n5120) );
  AND2_X1 U6284 ( .A1(n5239), .A2(n5659), .ZN(n5121) );
  INV_X1 U6285 ( .A(n5648), .ZN(n5645) );
  NAND2_X1 U6286 ( .A1(n7957), .A2(n9399), .ZN(n5648) );
  NAND2_X1 U6287 ( .A1(n6869), .A2(n6868), .ZN(n10480) );
  NOR2_X1 U6288 ( .A1(n9426), .A2(n5726), .ZN(n5122) );
  NOR2_X1 U6289 ( .A1(n7101), .A2(n7547), .ZN(n5123) );
  AND2_X1 U6290 ( .A1(n7321), .A2(n6481), .ZN(n5124) );
  NAND2_X1 U6291 ( .A1(n9334), .A2(n9588), .ZN(n5125) );
  AND2_X1 U6292 ( .A1(n9589), .A2(n9756), .ZN(n5126) );
  AND2_X1 U6293 ( .A1(n6488), .A2(n5638), .ZN(n5127) );
  INV_X1 U6294 ( .A(n6459), .ZN(n5351) );
  NOR2_X1 U6295 ( .A1(n9510), .A2(n9509), .ZN(n5128) );
  INV_X1 U6296 ( .A(n10525), .ZN(n10376) );
  NAND2_X1 U6297 ( .A1(n6626), .A2(n6625), .ZN(n10525) );
  INV_X1 U6298 ( .A(n10255), .ZN(n10975) );
  NAND2_X1 U6299 ( .A1(n6842), .A2(n6841), .ZN(n10255) );
  AND2_X1 U6300 ( .A1(n8821), .A2(n8819), .ZN(n5129) );
  INV_X1 U6301 ( .A(n9973), .ZN(n5431) );
  AND2_X1 U6302 ( .A1(n9321), .A2(n9389), .ZN(n5130) );
  AND2_X1 U6303 ( .A1(n5620), .A2(n8813), .ZN(n5131) );
  NAND2_X1 U6304 ( .A1(n9402), .A2(n8401), .ZN(n7199) );
  INV_X1 U6305 ( .A(n7199), .ZN(n5486) );
  AND2_X1 U6306 ( .A1(n5429), .A2(n5243), .ZN(n5132) );
  AND2_X1 U6307 ( .A1(n9802), .A2(n5255), .ZN(n5133) );
  NOR2_X1 U6308 ( .A1(n8811), .A2(n9666), .ZN(n5134) );
  NOR2_X1 U6309 ( .A1(n9853), .A2(n9852), .ZN(n5135) );
  NOR2_X1 U6310 ( .A1(n9806), .A2(n9805), .ZN(n5136) );
  NOR2_X1 U6311 ( .A1(n9657), .A2(n9669), .ZN(n5137) );
  NOR2_X1 U6312 ( .A1(n8619), .A2(n8609), .ZN(n5138) );
  AND2_X1 U6313 ( .A1(n8706), .A2(n9392), .ZN(n5139) );
  AND2_X1 U6314 ( .A1(n5564), .A2(n9501), .ZN(n5140) );
  INV_X1 U6315 ( .A(n5642), .ZN(n5641) );
  AND2_X1 U6316 ( .A1(n8303), .A2(n10881), .ZN(n5141) );
  INV_X1 U6317 ( .A(n5556), .ZN(n5555) );
  OAI21_X1 U6318 ( .B1(n5559), .B2(n5557), .A(n7335), .ZN(n5556) );
  INV_X1 U6319 ( .A(n5737), .ZN(n5670) );
  NOR2_X1 U6320 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5737) );
  AND2_X1 U6321 ( .A1(n5985), .A2(SI_7_), .ZN(n5142) );
  AND2_X1 U6322 ( .A1(n9760), .A2(n9602), .ZN(n5143) );
  AND2_X1 U6323 ( .A1(n6004), .A2(SI_12_), .ZN(n5144) );
  INV_X1 U6324 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5951) );
  OR2_X1 U6325 ( .A1(n5224), .A2(n9396), .ZN(n5145) );
  INV_X1 U6326 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9237) );
  AND2_X1 U6327 ( .A1(n8569), .A2(n8568), .ZN(n5146) );
  XNOR2_X1 U6328 ( .A(n6540), .B(n6541), .ZN(n7507) );
  NAND2_X1 U6329 ( .A1(n5807), .A2(n5734), .ZN(n5798) );
  AND2_X1 U6330 ( .A1(n7268), .A2(n7267), .ZN(n9659) );
  INV_X1 U6331 ( .A(n9659), .ZN(n5554) );
  NAND2_X1 U6332 ( .A1(n7107), .A2(n7021), .ZN(n5147) );
  AND2_X1 U6333 ( .A1(n7042), .A2(n10348), .ZN(n10362) );
  NAND2_X1 U6334 ( .A1(n7303), .A2(n7322), .ZN(n7348) );
  INV_X1 U6335 ( .A(n7348), .ZN(n5384) );
  AND2_X1 U6336 ( .A1(n6538), .A2(n6539), .ZN(n5148) );
  AND2_X1 U6337 ( .A1(n5552), .A2(n5112), .ZN(n5149) );
  AND2_X1 U6338 ( .A1(n5391), .A2(n5390), .ZN(n5150) );
  AND2_X1 U6339 ( .A1(n10447), .A2(n6888), .ZN(n5151) );
  AND2_X1 U6340 ( .A1(n5125), .A2(n7167), .ZN(n5152) );
  AND2_X1 U6341 ( .A1(n7299), .A2(n5301), .ZN(n5153) );
  AND2_X1 U6342 ( .A1(n7018), .A2(n7016), .ZN(n10548) );
  AND2_X1 U6343 ( .A1(n7782), .A2(n7781), .ZN(n5154) );
  OR2_X1 U6344 ( .A1(n7462), .A2(n10698), .ZN(n5155) );
  AND2_X1 U6345 ( .A1(n5362), .A2(n8529), .ZN(n5156) );
  AND2_X1 U6346 ( .A1(n7369), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5157) );
  AND2_X1 U6347 ( .A1(n5343), .A2(n5342), .ZN(n5158) );
  NAND2_X1 U6348 ( .A1(n9401), .A2(n7772), .ZN(n5159) );
  NAND2_X1 U6349 ( .A1(n7369), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5160) );
  AND2_X1 U6350 ( .A1(n5434), .A2(n9973), .ZN(n5161) );
  AND2_X1 U6351 ( .A1(n5113), .A2(n5741), .ZN(n5162) );
  AND2_X1 U6352 ( .A1(n5724), .A2(n5725), .ZN(n5163) );
  OR2_X1 U6353 ( .A1(n5816), .A2(n7641), .ZN(n5164) );
  AND2_X1 U6354 ( .A1(n5575), .A2(n5574), .ZN(n5165) );
  INV_X1 U6355 ( .A(n5717), .ZN(n5631) );
  INV_X1 U6356 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5778) );
  NOR2_X1 U6357 ( .A1(n9996), .A2(n5715), .ZN(n5166) );
  AND2_X1 U6358 ( .A1(n8837), .A2(n9386), .ZN(n5167) );
  AND4_X1 U6359 ( .A1(n6356), .A2(n6355), .A3(n6354), .A4(n6353), .ZN(n9654)
         );
  INV_X1 U6360 ( .A(n9654), .ZN(n5193) );
  INV_X1 U6361 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5427) );
  OAI21_X1 U6362 ( .B1(n8085), .B2(n6205), .A(n7218), .ZN(n8100) );
  OAI21_X1 U6363 ( .B1(n5751), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U6364 ( .A1(n5365), .A2(n5368), .ZN(n8460) );
  AND2_X1 U6365 ( .A1(n8644), .A2(n5399), .ZN(n5168) );
  NOR2_X1 U6366 ( .A1(n5108), .A2(n6689), .ZN(n6824) );
  OAI21_X1 U6367 ( .B1(n5222), .B2(n5221), .A(n5219), .ZN(n8763) );
  NAND2_X1 U6368 ( .A1(n8742), .A2(n8741), .ZN(n9803) );
  INV_X1 U6369 ( .A(n7739), .ZN(n7306) );
  NAND2_X1 U6370 ( .A1(n5194), .A2(n5553), .ZN(n9633) );
  INV_X1 U6371 ( .A(n5217), .ZN(n8664) );
  NAND2_X1 U6372 ( .A1(n8605), .A2(n8604), .ZN(n8739) );
  NAND2_X1 U6373 ( .A1(n5439), .A2(n8333), .ZN(n8566) );
  NAND2_X1 U6374 ( .A1(n5464), .A2(n5465), .ZN(n9658) );
  NAND2_X1 U6375 ( .A1(n5675), .A2(n8428), .ZN(n8556) );
  NAND2_X1 U6376 ( .A1(n6537), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6867) );
  NAND2_X1 U6377 ( .A1(n6950), .A2(n6949), .ZN(n10501) );
  INV_X1 U6378 ( .A(n10501), .ZN(n5414) );
  AND2_X1 U6379 ( .A1(n7706), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U6380 ( .A1(n5352), .A2(n6458), .ZN(n8722) );
  NOR2_X1 U6381 ( .A1(n6689), .A2(n6535), .ZN(n6822) );
  NOR2_X1 U6382 ( .A1(n8495), .A2(n5885), .ZN(n5170) );
  NAND2_X1 U6383 ( .A1(n10393), .A2(n5393), .ZN(n5394) );
  AND2_X1 U6384 ( .A1(n7873), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5171) );
  NAND2_X1 U6385 ( .A1(n9825), .A2(n9824), .ZN(n5172) );
  AND2_X1 U6386 ( .A1(n5887), .A2(n5495), .ZN(n5173) );
  AND2_X1 U6387 ( .A1(n9663), .A2(n5093), .ZN(n5174) );
  NAND2_X1 U6388 ( .A1(n7392), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5175) );
  AND2_X1 U6389 ( .A1(n5887), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5176) );
  INV_X1 U6390 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6536) );
  AND2_X1 U6391 ( .A1(n5630), .A2(n5629), .ZN(n5177) );
  INV_X1 U6392 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U6393 ( .A1(n9823), .A2(n10080), .ZN(n5178) );
  INV_X1 U6394 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9009) );
  NAND2_X1 U6395 ( .A1(n7949), .A2(n10472), .ZN(n10475) );
  INV_X2 U6396 ( .A(n10475), .ZN(n11005) );
  AND4_X1 U6397 ( .A1(n6622), .A2(n6621), .A3(n6620), .A4(n6619), .ZN(n10262)
         );
  INV_X1 U6398 ( .A(n10262), .ZN(n5699) );
  NAND2_X1 U6399 ( .A1(n6487), .A2(n6488), .ZN(n6490) );
  NAND2_X1 U6400 ( .A1(n7758), .A2(n7759), .ZN(n7757) );
  NAND2_X1 U6401 ( .A1(n8794), .A2(n7805), .ZN(n7825) );
  NAND2_X1 U6402 ( .A1(n5202), .A2(n5555), .ZN(n8265) );
  NAND2_X1 U6403 ( .A1(n8446), .A2(n8445), .ZN(n5179) );
  NAND2_X1 U6404 ( .A1(n5500), .A2(n7224), .ZN(n8085) );
  NAND2_X1 U6405 ( .A1(n5681), .A2(n8274), .ZN(n10877) );
  INV_X1 U6406 ( .A(n6465), .ZN(n6481) );
  NAND2_X1 U6407 ( .A1(n6880), .A2(n6879), .ZN(n10543) );
  INV_X1 U6408 ( .A(n10543), .ZN(n5396) );
  INV_X1 U6409 ( .A(n8528), .ZN(n5366) );
  NOR3_X1 U6410 ( .A1(n9720), .A2(n7739), .A3(P2_U3151), .ZN(n5180) );
  OAI21_X1 U6411 ( .B1(n5356), .B2(n5355), .A(n5353), .ZN(n7915) );
  INV_X1 U6412 ( .A(n10939), .ZN(n5526) );
  AND2_X1 U6413 ( .A1(n7176), .A2(n8528), .ZN(n8461) );
  NOR2_X1 U6414 ( .A1(n8208), .A2(n8207), .ZN(n5181) );
  INV_X1 U6415 ( .A(n5635), .ZN(n5634) );
  AND2_X1 U6416 ( .A1(n8666), .A2(n5117), .ZN(n5635) );
  INV_X1 U6417 ( .A(n5270), .ZN(n5269) );
  NOR2_X1 U6418 ( .A1(n6547), .A2(n9044), .ZN(n5270) );
  OR2_X1 U6419 ( .A1(n9489), .A2(n9468), .ZN(n5182) );
  INV_X1 U6420 ( .A(n5406), .ZN(n10947) );
  NOR2_X1 U6421 ( .A1(n10879), .A2(n5408), .ZN(n5406) );
  NOR3_X1 U6422 ( .A1(n10879), .A2(n10957), .A3(n5408), .ZN(n5405) );
  AND2_X1 U6423 ( .A1(n5214), .A2(n5154), .ZN(n7956) );
  AND2_X1 U6424 ( .A1(n6057), .A2(SI_25_), .ZN(n5183) );
  INV_X1 U6425 ( .A(n9445), .ZN(n5497) );
  XNOR2_X1 U6426 ( .A(n6555), .B(n9021), .ZN(n7151) );
  INV_X1 U6427 ( .A(n7991), .ZN(n7969) );
  XNOR2_X1 U6428 ( .A(n5786), .B(P2_IR_REG_19__SCAN_IN), .ZN(n6480) );
  AND2_X1 U6429 ( .A1(n6547), .A2(n9044), .ZN(n5184) );
  AND4_X1 U6430 ( .A1(n6860), .A2(n6859), .A3(n6858), .A4(n6857), .ZN(n10465)
         );
  INV_X1 U6431 ( .A(n10465), .ZN(n5693) );
  NAND2_X1 U6432 ( .A1(n6114), .A2(n6113), .ZN(n7666) );
  OR2_X1 U6433 ( .A1(n8047), .A2(n9397), .ZN(n5185) );
  INV_X1 U6434 ( .A(n7730), .ZN(n8122) );
  INV_X1 U6435 ( .A(n7508), .ZN(n5453) );
  NOR2_X1 U6436 ( .A1(n6481), .A2(n8122), .ZN(n5186) );
  NAND2_X1 U6437 ( .A1(n7698), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5187) );
  INV_X1 U6438 ( .A(n6480), .ZN(n8042) );
  XOR2_X1 U6439 ( .A(n10182), .B(P1_REG2_REG_16__SCAN_IN), .Z(n5188) );
  AND2_X1 U6440 ( .A1(n5479), .A2(n5478), .ZN(n5189) );
  INV_X1 U6441 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U6442 ( .A1(n5885), .A2(n5491), .ZN(n5489) );
  XNOR2_X1 U6443 ( .A(n5840), .B(n8505), .ZN(n8500) );
  NAND3_X1 U6444 ( .A1(n7144), .A2(n7140), .A3(n7546), .ZN(n7141) );
  INV_X1 U6445 ( .A(n7145), .ZN(n7166) );
  NAND2_X1 U6446 ( .A1(n10736), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5598) );
  INV_X1 U6447 ( .A(n6083), .ZN(n5594) );
  OAI21_X1 U6448 ( .B1(n6938), .B2(n7547), .A(n7041), .ZN(n5341) );
  INV_X1 U6449 ( .A(n5338), .ZN(n6964) );
  NAND2_X1 U6450 ( .A1(n5328), .A2(n5151), .ZN(n6911) );
  NAND2_X1 U6451 ( .A1(n6911), .A2(n5327), .ZN(n6908) );
  NAND2_X1 U6452 ( .A1(n6922), .A2(n6976), .ZN(n5337) );
  AOI22_X2 U6453 ( .A1(n10341), .A2(n10342), .B1(n10363), .B2(n10514), .ZN(
        n10329) );
  XNOR2_X2 U6454 ( .A(n7077), .B(n10776), .ZN(n7991) );
  NAND2_X2 U6455 ( .A1(n9547), .A2(n6483), .ZN(n6517) );
  AND2_X2 U6457 ( .A1(n5668), .A2(n5669), .ZN(n5776) );
  INV_X1 U6458 ( .A(n7767), .ZN(n5664) );
  INV_X1 U6459 ( .A(n5211), .ZN(n5210) );
  XNOR2_X1 U6460 ( .A(n7735), .B(n8312), .ZN(n5211) );
  NAND2_X1 U6461 ( .A1(n5215), .A2(n5162), .ZN(n5742) );
  CLKBUF_X1 U6462 ( .A(n5222), .Z(n5217) );
  AND2_X1 U6463 ( .A1(n5799), .A2(n5734), .ZN(n5227) );
  NAND4_X1 U6464 ( .A1(n5807), .A2(n5227), .A3(n5228), .A4(n5083), .ZN(n5791)
         );
  NAND2_X1 U6465 ( .A1(n9372), .A2(n5232), .ZN(n5231) );
  OAI211_X1 U6466 ( .C1(n9372), .C2(n5233), .A(n5231), .B(n9285), .ZN(P2_U3160) );
  NAND2_X1 U6467 ( .A1(n5241), .A2(n5582), .ZN(n5240) );
  NAND2_X1 U6468 ( .A1(n5977), .A2(n5581), .ZN(n5241) );
  NAND2_X1 U6469 ( .A1(n6122), .A2(n6123), .ZN(n5977) );
  NAND2_X1 U6470 ( .A1(n5428), .A2(n5429), .ZN(n9865) );
  NAND2_X1 U6471 ( .A1(n10048), .A2(n10049), .ZN(n5242) );
  INV_X1 U6472 ( .A(n9864), .ZN(n5243) );
  NAND2_X1 U6473 ( .A1(n6207), .A2(n5614), .ZN(n5250) );
  OAI21_X1 U6474 ( .B1(n6207), .B2(n5249), .A(n5247), .ZN(n6245) );
  NAND2_X1 U6475 ( .A1(n5246), .A2(n5245), .ZN(n6007) );
  AOI21_X1 U6476 ( .B1(n5247), .B2(n5249), .A(n6244), .ZN(n5246) );
  NAND3_X1 U6477 ( .A1(n8605), .A2(n5256), .A3(n8604), .ZN(n5253) );
  NAND3_X1 U6478 ( .A1(n8605), .A2(n8604), .A3(n5711), .ZN(n5254) );
  INV_X1 U6479 ( .A(n8744), .ZN(n8742) );
  NAND2_X1 U6480 ( .A1(n6067), .A2(n5107), .ZN(n5258) );
  NAND2_X1 U6481 ( .A1(n6067), .A2(n6051), .ZN(n6374) );
  INV_X2 U6482 ( .A(n9953), .ZN(n9901) );
  NAND3_X1 U6483 ( .A1(n5276), .A2(n5273), .A3(n5371), .ZN(n5374) );
  NAND3_X1 U6484 ( .A1(n5275), .A2(n5599), .A3(n5274), .ZN(n5273) );
  NAND2_X1 U6485 ( .A1(n9983), .A2(n9984), .ZN(n9982) );
  NAND2_X1 U6486 ( .A1(n9982), .A2(n9892), .ZN(n10069) );
  AND3_X2 U6487 ( .A1(n5163), .A2(n5682), .A3(n5283), .ZN(n6988) );
  NOR2_X2 U6488 ( .A1(n6535), .A2(n5683), .ZN(n5682) );
  NAND3_X1 U6489 ( .A1(n7330), .A2(n5286), .A3(n5285), .ZN(n5284) );
  NAND2_X1 U6490 ( .A1(n5965), .A2(n5288), .ZN(n5968) );
  NAND3_X1 U6491 ( .A1(n5597), .A2(n5595), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n5288) );
  INV_X2 U6492 ( .A(n5974), .ZN(n7361) );
  AOI21_X1 U6493 ( .B1(n9511), .B2(n9513), .A(n5290), .ZN(n5863) );
  INV_X2 U6494 ( .A(n5813), .ZN(n5871) );
  NOR2_X1 U6495 ( .A1(n9566), .A2(n7293), .ZN(n5300) );
  OAI211_X1 U6496 ( .C1(n7294), .C2(n5296), .A(n5384), .B(n5294), .ZN(n5303)
         );
  AOI21_X1 U6497 ( .B1(n5295), .B2(n7300), .A(n5303), .ZN(n7307) );
  OAI21_X1 U6498 ( .B1(n5305), .B2(n8126), .A(n5304), .ZN(n5840) );
  OAI21_X1 U6499 ( .B1(n7441), .B2(n5308), .A(n5307), .ZN(n7483) );
  NAND2_X1 U6500 ( .A1(n5911), .A2(n5309), .ZN(n5308) );
  NOR2_X1 U6501 ( .A1(n7441), .A2(n5819), .ZN(n5820) );
  NOR2_X1 U6502 ( .A1(n7483), .A2(n8400), .ZN(n7482) );
  NAND3_X1 U6503 ( .A1(n5312), .A2(n7251), .A3(n7253), .ZN(n5311) );
  NAND3_X1 U6504 ( .A1(n7248), .A2(n7250), .A3(n7249), .ZN(n5312) );
  INV_X1 U6505 ( .A(n6452), .ZN(n5315) );
  NAND2_X1 U6506 ( .A1(n5316), .A2(n5313), .ZN(n7239) );
  NOR2_X1 U6507 ( .A1(n5315), .A2(n7306), .ZN(n5314) );
  NAND3_X1 U6508 ( .A1(n5323), .A2(n5320), .A3(n5319), .ZN(n5318) );
  NAND3_X1 U6509 ( .A1(n7259), .A2(n7257), .A3(n5321), .ZN(n5320) );
  NAND4_X1 U6510 ( .A1(n7266), .A2(n7263), .A3(n7265), .A4(n5324), .ZN(n5323)
         );
  INV_X4 U6511 ( .A(n7361), .ZN(n7362) );
  MUX2_X1 U6512 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7361), .Z(n5985) );
  NAND3_X1 U6513 ( .A1(n5326), .A2(n5325), .A3(n5989), .ZN(n6194) );
  NAND3_X1 U6514 ( .A1(n5585), .A2(n5584), .A3(n6174), .ZN(n5325) );
  NAND3_X1 U6515 ( .A1(n5585), .A2(n5584), .A3(n5983), .ZN(n5326) );
  NAND3_X1 U6516 ( .A1(n5331), .A2(n5330), .A3(n5329), .ZN(n5328) );
  NAND3_X1 U6517 ( .A1(n6756), .A2(n6755), .A3(n5158), .ZN(n6786) );
  NAND3_X1 U6518 ( .A1(n6747), .A2(n8186), .A3(n6748), .ZN(n5342) );
  NAND4_X1 U6519 ( .A1(n6754), .A2(n6753), .A3(n8186), .A4(n6752), .ZN(n5343)
         );
  MUX2_X1 U6520 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7361), .Z(n5979) );
  INV_X1 U6521 ( .A(n5978), .ZN(n5345) );
  MUX2_X1 U6522 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n7361), .Z(n5346) );
  NAND2_X1 U6523 ( .A1(n5347), .A2(n5115), .ZN(n6087) );
  INV_X1 U6524 ( .A(n6162), .ZN(n5347) );
  NAND2_X1 U6525 ( .A1(n6475), .A2(n7362), .ZN(n6162) );
  OAI21_X1 U6526 ( .B1(n7759), .B2(n5357), .A(n7920), .ZN(n5354) );
  OR2_X1 U6527 ( .A1(n5357), .A2(n5358), .ZN(n5356) );
  NAND2_X1 U6528 ( .A1(n9626), .A2(n5360), .ZN(n5359) );
  NAND2_X1 U6529 ( .A1(n5359), .A2(n5152), .ZN(n6461) );
  NAND2_X1 U6530 ( .A1(n8268), .A2(n5364), .ZN(n5363) );
  NAND2_X1 U6531 ( .A1(n5363), .A2(n5156), .ZN(n8530) );
  NAND2_X1 U6532 ( .A1(n5374), .A2(n7357), .ZN(P2_U3296) );
  NAND2_X1 U6533 ( .A1(n9696), .A2(n5385), .ZN(n5388) );
  NAND2_X1 U6534 ( .A1(n5376), .A2(n5380), .ZN(n7324) );
  NAND2_X1 U6535 ( .A1(n9696), .A2(n5377), .ZN(n5376) );
  NAND2_X1 U6536 ( .A1(n5388), .A2(n7292), .ZN(n9557) );
  OAI21_X2 U6537 ( .B1(n5379), .B2(n5387), .A(n6463), .ZN(n7323) );
  NOR2_X2 U6538 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6664) );
  NAND2_X1 U6539 ( .A1(n6664), .A2(n5389), .ZN(n6687) );
  INV_X1 U6540 ( .A(n5394), .ZN(n10357) );
  NAND2_X1 U6541 ( .A1(n6988), .A2(n5401), .ZN(n5404) );
  INV_X1 U6542 ( .A(n5405), .ZN(n10948) );
  NOR2_X1 U6543 ( .A1(n10320), .A2(n5412), .ZN(n10275) );
  NOR2_X1 U6544 ( .A1(n10320), .A2(n10501), .ZN(n10307) );
  AND2_X2 U6545 ( .A1(n6649), .A2(n5415), .ZN(n10776) );
  NAND2_X1 U6546 ( .A1(n5419), .A2(n5188), .ZN(n10181) );
  OR2_X1 U6547 ( .A1(n10168), .A2(n10169), .ZN(n5419) );
  NAND2_X1 U6548 ( .A1(n9937), .A2(n5161), .ZN(n5428) );
  NAND2_X1 U6549 ( .A1(n8329), .A2(n5440), .ZN(n5437) );
  NAND2_X1 U6550 ( .A1(n5437), .A2(n5438), .ZN(n8575) );
  NAND2_X1 U6551 ( .A1(n5445), .A2(n5166), .ZN(n5444) );
  INV_X1 U6552 ( .A(n5445), .ZN(n9995) );
  NAND2_X1 U6553 ( .A1(n5444), .A2(n5172), .ZN(n10005) );
  INV_X1 U6554 ( .A(n7829), .ZN(n5448) );
  NAND2_X1 U6555 ( .A1(n8146), .A2(n8145), .ZN(n5449) );
  NAND2_X1 U6556 ( .A1(n8156), .A2(n8157), .ZN(n8299) );
  NAND3_X1 U6557 ( .A1(n5449), .A2(n8147), .A3(n8161), .ZN(n8156) );
  NAND2_X1 U6558 ( .A1(n6867), .A2(n5148), .ZN(n6893) );
  NAND2_X2 U6559 ( .A1(n5454), .A2(n7511), .ZN(n9860) );
  NAND2_X2 U6560 ( .A1(n7510), .A2(n7511), .ZN(n9951) );
  NAND2_X1 U6561 ( .A1(n8070), .A2(n8069), .ZN(n8146) );
  XNOR2_X2 U6562 ( .A(n5457), .B(P2_IR_REG_1__SCAN_IN), .ZN(n5868) );
  INV_X1 U6563 ( .A(n5460), .ZN(n9480) );
  INV_X1 U6564 ( .A(n5458), .ZN(n9478) );
  NOR2_X1 U6565 ( .A1(n9461), .A2(n9462), .ZN(n9460) );
  NAND2_X1 U6566 ( .A1(n6460), .A2(n5099), .ZN(n5463) );
  NAND2_X1 U6567 ( .A1(n6460), .A2(n7260), .ZN(n9675) );
  INV_X1 U6568 ( .A(n7265), .ZN(n5468) );
  OAI211_X1 U6569 ( .C1(n5817), .C2(n7641), .A(n5469), .B(n5164), .ZN(n7439)
         );
  NAND3_X1 U6570 ( .A1(n5816), .A2(n5817), .A3(n7641), .ZN(n5469) );
  NAND2_X1 U6571 ( .A1(n5870), .A2(n5470), .ZN(n5473) );
  INV_X1 U6572 ( .A(n5479), .ZN(n7478) );
  INV_X1 U6573 ( .A(n5874), .ZN(n5478) );
  OR2_X2 U6574 ( .A1(n10715), .A2(n5483), .ZN(n5482) );
  INV_X1 U6575 ( .A(n5485), .ZN(n10714) );
  INV_X1 U6576 ( .A(n5878), .ZN(n5484) );
  NAND2_X1 U6577 ( .A1(n7681), .A2(n7682), .ZN(n7680) );
  OAI21_X1 U6578 ( .B1(n8496), .B2(n5490), .A(n5489), .ZN(n9416) );
  NAND2_X1 U6579 ( .A1(n5889), .A2(n5497), .ZN(n5493) );
  NAND2_X1 U6580 ( .A1(n5493), .A2(n5492), .ZN(n9444) );
  NAND3_X1 U6581 ( .A1(n5496), .A2(n5887), .A3(n5494), .ZN(n5492) );
  OR2_X2 U6582 ( .A1(n5888), .A2(n7472), .ZN(n5496) );
  NAND2_X1 U6583 ( .A1(n5496), .A2(n5887), .ZN(n9438) );
  NAND2_X2 U6584 ( .A1(n6453), .A2(n7237), .ZN(n8268) );
  NAND2_X1 U6585 ( .A1(n5776), .A2(n5774), .ZN(n5779) );
  CLKBUF_X1 U6586 ( .A(n5776), .Z(n5501) );
  XNOR2_X1 U6587 ( .A(n7323), .B(n7348), .ZN(n9545) );
  NOR2_X2 U6588 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5503) );
  NOR2_X1 U6589 ( .A1(n8020), .A2(n7991), .ZN(n7050) );
  INV_X1 U6590 ( .A(n8550), .ZN(n5506) );
  NAND2_X1 U6591 ( .A1(n5506), .A2(n7058), .ZN(n5508) );
  NAND2_X1 U6592 ( .A1(n5508), .A2(n5507), .ZN(n7019) );
  AND2_X1 U6593 ( .A1(n10548), .A2(n5509), .ZN(n5507) );
  OAI22_X2 U6594 ( .A1(n10377), .A2(n5512), .B1(n5513), .B2(n10240), .ZN(
        n10335) );
  NAND2_X1 U6595 ( .A1(n10335), .A2(n10334), .ZN(n10333) );
  NAND2_X1 U6596 ( .A1(n6560), .A2(n9236), .ZN(n6562) );
  NOR2_X1 U6597 ( .A1(n10303), .A2(n10302), .ZN(n10301) );
  OAI21_X2 U6598 ( .B1(n10459), .B2(n5147), .A(n5529), .ZN(n10432) );
  OAI21_X1 U6599 ( .B1(n8012), .B2(n5534), .A(n5533), .ZN(n8184) );
  OAI21_X1 U6600 ( .B1(n8012), .B2(n7003), .A(n7088), .ZN(n7988) );
  OAI21_X1 U6601 ( .B1(n8458), .B2(n5541), .A(n5538), .ZN(n6281) );
  NAND2_X1 U6602 ( .A1(n6294), .A2(n5546), .ZN(n5544) );
  NAND2_X1 U6603 ( .A1(n6294), .A2(n6293), .ZN(n8720) );
  NAND2_X1 U6604 ( .A1(n5776), .A2(n5561), .ZN(n5953) );
  NAND2_X1 U6605 ( .A1(n5776), .A2(n5106), .ZN(n9781) );
  NAND2_X1 U6606 ( .A1(n9424), .A2(n5567), .ZN(n5565) );
  NAND2_X1 U6607 ( .A1(n5566), .A2(n5565), .ZN(n9450) );
  INV_X1 U6608 ( .A(n5850), .ZN(n5574) );
  NAND2_X1 U6609 ( .A1(n5850), .A2(n5573), .ZN(n5572) );
  INV_X1 U6610 ( .A(n5575), .ZN(n9467) );
  INV_X1 U6611 ( .A(n5580), .ZN(n5582) );
  NAND2_X1 U6612 ( .A1(n5583), .A2(n5978), .ZN(n6147) );
  NAND2_X1 U6613 ( .A1(n6136), .A2(n6137), .ZN(n5583) );
  NAND2_X1 U6614 ( .A1(n6657), .A2(n6096), .ZN(n6083) );
  INV_X1 U6615 ( .A(n7305), .ZN(n5604) );
  AOI21_X1 U6616 ( .B1(n7307), .B2(n7306), .A(n7326), .ZN(n5603) );
  NAND2_X1 U6617 ( .A1(n6256), .A2(n5612), .ZN(n5608) );
  OAI21_X1 U6618 ( .B1(n6256), .B2(n6255), .A(n6011), .ZN(n6268) );
  XNOR2_X1 U6619 ( .A(n7734), .B(n5619), .ZN(n7936) );
  INV_X1 U6620 ( .A(n9404), .ZN(n5619) );
  NAND2_X1 U6621 ( .A1(n7934), .A2(n5119), .ZN(n7927) );
  INV_X1 U6622 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5638) );
  INV_X1 U6623 ( .A(n7956), .ZN(n5644) );
  NOR2_X1 U6624 ( .A1(n7956), .A2(n5645), .ZN(n7958) );
  INV_X1 U6625 ( .A(n9398), .ZN(n5647) );
  NAND2_X1 U6626 ( .A1(n9372), .A2(n5650), .ZN(n5649) );
  OAI211_X1 U6627 ( .C1(n9372), .C2(n5651), .A(n5649), .B(n8842), .ZN(n5657)
         );
  XNOR2_X1 U6628 ( .A(n5657), .B(n9254), .ZN(P2_U3154) );
  INV_X1 U6629 ( .A(n9279), .ZN(n5659) );
  NAND3_X1 U6630 ( .A1(n7742), .A2(n5666), .A3(n7777), .ZN(n5663) );
  NAND2_X1 U6631 ( .A1(n9262), .A2(n5667), .ZN(n9295) );
  NAND3_X1 U6632 ( .A1(n5668), .A2(n5669), .A3(n5761), .ZN(n5753) );
  NAND2_X1 U6633 ( .A1(n5671), .A2(n5673), .ZN(n10937) );
  NAND2_X1 U6634 ( .A1(n8426), .A2(n5672), .ZN(n5671) );
  NAND2_X1 U6635 ( .A1(n5676), .A2(n5678), .ZN(n8371) );
  NAND2_X1 U6636 ( .A1(n8273), .A2(n5677), .ZN(n5676) );
  NAND2_X1 U6637 ( .A1(n5283), .A2(n5682), .ZN(n6542) );
  NAND2_X2 U6638 ( .A1(n10314), .A2(n10315), .ZN(n10313) );
  NAND2_X1 U6639 ( .A1(n10547), .A2(n5689), .ZN(n5686) );
  NAND2_X1 U6640 ( .A1(n5686), .A2(n5687), .ZN(n10446) );
  CLKBUF_X1 U6641 ( .A(n5696), .Z(n5694) );
  NAND2_X1 U6642 ( .A1(n10421), .A2(n5718), .ZN(n10401) );
  INV_X1 U6643 ( .A(n5718), .ZN(n5698) );
  AND2_X1 U6644 ( .A1(n6554), .A2(n5703), .ZN(n7155) );
  NAND2_X1 U6645 ( .A1(n6554), .A2(n5701), .ZN(n5700) );
  NAND2_X1 U6646 ( .A1(n6554), .A2(n6553), .ZN(n7158) );
  NAND2_X1 U6647 ( .A1(n6449), .A2(n6448), .ZN(n7671) );
  INV_X1 U6648 ( .A(n6064), .ZN(n6066) );
  INV_X1 U6649 ( .A(n8575), .ZN(n8573) );
  XNOR2_X1 U6650 ( .A(n5771), .B(n5772), .ZN(n7721) );
  NAND2_X1 U6651 ( .A1(n6393), .A2(n9387), .ZN(n6394) );
  XNOR2_X1 U6652 ( .A(n6549), .B(SI_29_), .ZN(n8789) );
  INV_X1 U6653 ( .A(n7495), .ZN(n8780) );
  NAND2_X1 U6654 ( .A1(n7494), .A2(n7495), .ZN(n10574) );
  INV_X1 U6655 ( .A(n7327), .ZN(n7321) );
  NAND2_X1 U6656 ( .A1(n5974), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U6657 ( .A1(n9628), .A2(n9627), .ZN(n9626) );
  XNOR2_X1 U6658 ( .A(n6399), .B(n6398), .ZN(n8779) );
  NAND2_X1 U6659 ( .A1(n9595), .A2(n9594), .ZN(n9702) );
  INV_X1 U6660 ( .A(n10005), .ZN(n10010) );
  INV_X1 U6661 ( .A(n5956), .ZN(n9259) );
  NOR2_X2 U6662 ( .A1(n7646), .A2(n7645), .ZN(n7652) );
  NAND2_X1 U6663 ( .A1(n7657), .A2(n7797), .ZN(n7081) );
  INV_X1 U6664 ( .A(n7657), .ZN(n7812) );
  OR2_X1 U6665 ( .A1(n7155), .A2(n6838), .ZN(n7156) );
  NOR2_X1 U6666 ( .A1(n6199), .A2(n6183), .ZN(n5707) );
  INV_X1 U6667 ( .A(n8086), .ZN(n6205) );
  OR2_X1 U6668 ( .A1(n9368), .A2(n9602), .ZN(n5708) );
  XOR2_X1 U6669 ( .A(n9514), .B(n9513), .Z(n5709) );
  XOR2_X1 U6670 ( .A(n5939), .B(n5863), .Z(n5710) );
  NAND2_X1 U6671 ( .A1(n8610), .A2(n8611), .ZN(n5711) );
  OR2_X1 U6672 ( .A1(n8436), .A2(n8435), .ZN(n5712) );
  AND2_X1 U6673 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5713) );
  INV_X1 U6674 ( .A(n5911), .ZN(n7491) );
  INV_X1 U6675 ( .A(n10702), .ZN(n7371) );
  AND2_X1 U6676 ( .A1(n7698), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5714) );
  AND2_X2 U6677 ( .A1(n8358), .A2(n9590), .ZN(n9673) );
  INV_X1 U6678 ( .A(n9405), .ZN(n6447) );
  AND2_X1 U6679 ( .A1(n9998), .A2(n9997), .ZN(n5715) );
  OR2_X1 U6680 ( .A1(n11008), .A2(n10450), .ZN(n5716) );
  AND2_X1 U6681 ( .A1(n8810), .A2(n8809), .ZN(n5717) );
  INV_X1 U6682 ( .A(n7630), .ZN(n6482) );
  INV_X1 U6683 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8417) );
  AND2_X1 U6684 ( .A1(n9752), .A2(n9576), .ZN(n5723) );
  AND3_X1 U6685 ( .A1(n9211), .A2(n9217), .A3(n6541), .ZN(n5724) );
  AND2_X1 U6686 ( .A1(n9212), .A2(n6539), .ZN(n5725) );
  AND2_X1 U6687 ( .A1(n5846), .A2(n7472), .ZN(n5726) );
  INV_X1 U6688 ( .A(n10271), .ZN(n10306) );
  NAND2_X1 U6689 ( .A1(n10746), .A2(n7656), .ZN(n10464) );
  INV_X1 U6690 ( .A(n10464), .ZN(n10550) );
  AND2_X1 U6691 ( .A1(n5993), .A2(n5992), .ZN(n5727) );
  NAND2_X1 U6692 ( .A1(n7731), .A2(n6504), .ZN(n9664) );
  AND3_X1 U6693 ( .A1(n10273), .A2(n10283), .A3(n7069), .ZN(n5728) );
  OR2_X1 U6694 ( .A1(n10734), .A2(n9524), .ZN(n5729) );
  NOR2_X1 U6695 ( .A1(n9966), .A2(n10064), .ZN(n5730) );
  NOR2_X2 U6696 ( .A1(n6574), .A2(n8790), .ZN(n5731) );
  INV_X1 U6697 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9217) );
  NAND2_X1 U6698 ( .A1(n5859), .A2(n6297), .ZN(n5860) );
  INV_X1 U6699 ( .A(n7884), .ZN(n6451) );
  INV_X1 U6700 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6543) );
  INV_X1 U6701 ( .A(n8449), .ZN(n8252) );
  AND2_X1 U6702 ( .A1(n7363), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5819) );
  AND3_X1 U6703 ( .A1(n9226), .A2(n9009), .A3(n9221), .ZN(n6553) );
  INV_X1 U6704 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7848) );
  NOR2_X1 U6705 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5781) );
  INV_X1 U6706 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8114) );
  OAI22_X1 U6707 ( .A1(n7919), .A2(n6165), .B1(n9399), .B2(n7790), .ZN(n7885)
         );
  AND2_X1 U6708 ( .A1(n5739), .A2(n5738), .ZN(n5749) );
  INV_X1 U6709 ( .A(n10008), .ZN(n9829) );
  INV_X1 U6710 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6763) );
  NAND2_X1 U6711 ( .A1(n7976), .A2(n7647), .ZN(n7515) );
  AND2_X1 U6712 ( .A1(n6637), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6618) );
  OR2_X1 U6713 ( .A1(n6773), .A2(n6772), .ZN(n6775) );
  INV_X1 U6714 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9001) );
  INV_X1 U6715 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6533) );
  INV_X1 U6716 ( .A(n9326), .ZN(n8828) );
  INV_X1 U6717 ( .A(n9348), .ZN(n8821) );
  INV_X1 U6718 ( .A(n6115), .ZN(n6128) );
  XNOR2_X1 U6719 ( .A(n5873), .B(n5911), .ZN(n7479) );
  OAI22_X1 U6720 ( .A1(n10659), .A2(n9637), .B1(n9635), .B2(n9589), .ZN(n9563)
         );
  OR2_X1 U6721 ( .A1(n9401), .A2(n8312), .ZN(n7200) );
  INV_X1 U6722 ( .A(n6518), .ZN(n6505) );
  INV_X1 U6723 ( .A(n8745), .ZN(n8741) );
  OAI211_X1 U6724 ( .C1(n7950), .C2(n7137), .A(n7136), .B(n5100), .ZN(n7138)
         );
  OR2_X1 U6725 ( .A1(n6844), .A2(n6843), .ZN(n6855) );
  AND2_X1 U6726 ( .A1(n6791), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6812) );
  AND2_X1 U6727 ( .A1(n7509), .A2(n7161), .ZN(n7656) );
  AOI22_X1 U6728 ( .A1(n10437), .A2(n10261), .B1(n10451), .B2(n11020), .ZN(
        n10420) );
  INV_X1 U6729 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9021) );
  INV_X1 U6730 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9017) );
  INV_X1 U6731 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6539) );
  AND2_X1 U6732 ( .A1(n6349), .A2(n9289), .ZN(n6362) );
  INV_X1 U6733 ( .A(n9402), .ZN(n7770) );
  OR2_X1 U6734 ( .A1(n7748), .A2(n7747), .ZN(n9361) );
  INV_X1 U6735 ( .A(n9330), .ZN(n9376) );
  OR2_X1 U6736 ( .A1(n6102), .A2(n9332), .ZN(n6380) );
  OR2_X1 U6737 ( .A1(n6102), .A2(n6351), .ZN(n6354) );
  OR2_X1 U6738 ( .A1(n5086), .A2(n10664), .ZN(n6080) );
  INV_X1 U6739 ( .A(n9551), .ZN(n9552) );
  OR2_X1 U6740 ( .A1(n9735), .A2(n6440), .ZN(n6529) );
  NAND2_X1 U6741 ( .A1(n9545), .A2(n6482), .ZN(n6483) );
  INV_X1 U6742 ( .A(n9666), .ZN(n9316) );
  INV_X1 U6743 ( .A(n9664), .ZN(n9653) );
  OR2_X1 U6744 ( .A1(n6490), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6492) );
  NAND2_X1 U6745 ( .A1(n8573), .A2(n8572), .ZN(n8604) );
  NOR2_X1 U6746 ( .A1(n9872), .A2(n9871), .ZN(n10016) );
  OR2_X1 U6747 ( .A1(n6829), .A2(n6828), .ZN(n6844) );
  AND2_X1 U6748 ( .A1(n7528), .A2(n10573), .ZN(n7524) );
  INV_X1 U6749 ( .A(n8788), .ZN(n10746) );
  NAND2_X1 U6750 ( .A1(n5731), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6671) );
  AND2_X1 U6751 ( .A1(n8384), .A2(n8383), .ZN(n8387) );
  OR2_X1 U6752 ( .A1(n10163), .A2(n10164), .ZN(n10176) );
  AND2_X1 U6753 ( .A1(n5452), .A2(n8123), .ZN(n7540) );
  AND4_X1 U6754 ( .A1(n6947), .A2(n6946), .A3(n6945), .A4(n6944), .ZN(n10305)
         );
  INV_X1 U6755 ( .A(n10417), .ZN(n10451) );
  AND2_X1 U6756 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6720) );
  INV_X1 U6757 ( .A(n10260), .ZN(n11020) );
  INV_X1 U6758 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9226) );
  XNOR2_X1 U6759 ( .A(n6004), .B(n8869), .ZN(n6231) );
  INV_X1 U6760 ( .A(n9328), .ZN(n9380) );
  OR2_X1 U6761 ( .A1(n6102), .A2(n9533), .ZN(n7318) );
  AND4_X1 U6762 ( .A1(n6382), .A2(n6381), .A3(n6380), .A4(n6379), .ZN(n9588)
         );
  OR2_X1 U6763 ( .A1(n5085), .A2(n7480), .ZN(n6120) );
  NOR2_X1 U6764 ( .A1(n5876), .A2(n10693), .ZN(n7456) );
  NOR2_X1 U6765 ( .A1(n5881), .A2(n8136), .ZN(n8200) );
  AOI21_X1 U6766 ( .B1(n5946), .B2(n10729), .A(n5945), .ZN(n5947) );
  NAND2_X1 U6767 ( .A1(n8530), .A2(n6456), .ZN(n8624) );
  INV_X1 U6768 ( .A(n9590), .ZN(n10871) );
  AND2_X1 U6769 ( .A1(n10874), .A2(n10865), .ZN(n9677) );
  OAI21_X1 U6770 ( .B1(n9542), .B2(n9738), .A(n6529), .ZN(n6530) );
  AND2_X1 U6771 ( .A1(n6520), .A2(n6519), .ZN(n8242) );
  INV_X1 U6772 ( .A(n9733), .ZN(n9718) );
  OR2_X1 U6773 ( .A1(n8292), .A2(n6482), .ZN(n9733) );
  OAI21_X1 U6774 ( .B1(n7746), .B2(n6509), .A(n6508), .ZN(n6512) );
  AND2_X1 U6775 ( .A1(n5857), .A2(n5856), .ZN(n9493) );
  INV_X1 U6776 ( .A(n10041), .ZN(n10029) );
  AND4_X1 U6777 ( .A1(n6960), .A2(n6959), .A3(n6958), .A4(n6957), .ZN(n10319)
         );
  AND4_X1 U6778 ( .A1(n6632), .A2(n6631), .A3(n6630), .A4(n6629), .ZN(n10264)
         );
  AND4_X1 U6779 ( .A1(n6834), .A2(n6833), .A3(n6832), .A4(n6831), .ZN(n9924)
         );
  AND2_X1 U6780 ( .A1(n8222), .A2(n8221), .ZN(n10114) );
  INV_X1 U6781 ( .A(n10756), .ZN(n10203) );
  NOR2_X1 U6782 ( .A1(n7569), .A2(n7568), .ZN(n10222) );
  AND2_X1 U6783 ( .A1(n7540), .A2(n7525), .ZN(n10949) );
  NAND2_X1 U6784 ( .A1(n7041), .A2(n7040), .ZN(n10315) );
  NAND2_X1 U6785 ( .A1(n7975), .A2(n10997), .ZN(n10961) );
  AND2_X1 U6786 ( .A1(n7543), .A2(n7550), .ZN(n7944) );
  INV_X1 U6787 ( .A(n10848), .ZN(n10990) );
  NAND2_X1 U6788 ( .A1(n10848), .A2(n10928), .ZN(n11022) );
  AND2_X1 U6789 ( .A1(n6787), .A2(n6760), .ZN(n10105) );
  NAND2_X1 U6790 ( .A1(n7740), .A2(n5180), .ZN(n9355) );
  INV_X1 U6791 ( .A(n9364), .ZN(n9377) );
  AND4_X1 U6792 ( .A1(n7318), .A2(n6444), .A3(n6443), .A4(n6442), .ZN(n9550)
         );
  OR2_X1 U6793 ( .A1(P2_U3150), .A2(n5866), .ZN(n10734) );
  NAND2_X1 U6794 ( .A1(n7425), .A2(n7353), .ZN(n10724) );
  OAI21_X1 U6795 ( .B1(n5948), .B2(n10717), .A(n5947), .ZN(n5949) );
  INV_X1 U6796 ( .A(n6530), .ZN(n6531) );
  AND2_X2 U6797 ( .A1(n8242), .A2(n6528), .ZN(n9735) );
  AND3_X1 U6798 ( .A1(n8296), .A2(n8104), .A3(n8103), .ZN(n10923) );
  AND2_X2 U6799 ( .A1(n6512), .A2(n7397), .ZN(n11017) );
  NAND2_X1 U6800 ( .A1(n6512), .A2(n6511), .ZN(n9779) );
  AND2_X1 U6801 ( .A1(n7722), .A2(n8783), .ZN(n7397) );
  INV_X1 U6802 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8108) );
  INV_X1 U6803 ( .A(n9790), .ZN(n9783) );
  AND2_X1 U6804 ( .A1(n7413), .A2(n7412), .ZN(n10756) );
  INV_X1 U6805 ( .A(n10480), .ZN(n11008) );
  INV_X1 U6806 ( .A(n10071), .ZN(n10084) );
  INV_X1 U6807 ( .A(n10073), .ZN(n10090) );
  AND4_X1 U6808 ( .A1(n6584), .A2(n6583), .A3(n6582), .A4(n6581), .ZN(n9960)
         );
  AND4_X1 U6809 ( .A1(n6641), .A2(n6640), .A3(n6639), .A4(n6638), .ZN(n10433)
         );
  INV_X1 U6810 ( .A(n10959), .ZN(n10477) );
  INV_X1 U6811 ( .A(n10961), .ZN(n10458) );
  INV_X1 U6812 ( .A(n10475), .ZN(n10955) );
  INV_X1 U6813 ( .A(n11037), .ZN(n11035) );
  INV_X1 U6814 ( .A(n11041), .ZN(n11038) );
  AND2_X2 U6815 ( .A1(n7552), .A2(n7946), .ZN(n11041) );
  INV_X1 U6816 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n9155) );
  OR2_X1 U6817 ( .A1(n6840), .A2(n6839), .ZN(n10131) );
  INV_X1 U6818 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7418) );
  NAND2_X1 U6819 ( .A1(n6516), .A2(n6515), .ZN(P2_U3456) );
  INV_X2 U6820 ( .A(n10104), .ZN(P1_U3973) );
  NOR2_X1 U6821 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5739) );
  NOR2_X1 U6822 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5738) );
  INV_X1 U6823 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5741) );
  NAND2_X1 U6824 ( .A1(n5786), .A2(n5747), .ZN(n5743) );
  INV_X1 U6825 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U6826 ( .A1(n6446), .A2(n5744), .ZN(n5745) );
  NOR3_X1 U6827 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .A3(
        P2_IR_REG_13__SCAN_IN), .ZN(n5748) );
  NAND4_X1 U6828 ( .A1(n5749), .A2(n5748), .A3(n5747), .A4(n5741), .ZN(n5750)
         );
  NAND2_X1 U6829 ( .A1(n5771), .A2(n5772), .ZN(n5754) );
  NAND2_X1 U6830 ( .A1(n5759), .A2(n5758), .ZN(n5755) );
  INV_X1 U6831 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5756) );
  INV_X1 U6832 ( .A(n6485), .ZN(n5769) );
  INV_X1 U6833 ( .A(n6484), .ZN(n5767) );
  NOR3_X1 U6834 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5760) );
  NAND2_X1 U6835 ( .A1(n5762), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5763) );
  MUX2_X1 U6836 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5763), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5766) );
  INV_X1 U6837 ( .A(n7722), .ZN(n5770) );
  OR2_X1 U6838 ( .A1(n7739), .A2(n5770), .ZN(n5773) );
  NAND2_X1 U6839 ( .A1(n5773), .A2(n7721), .ZN(n5943) );
  NAND2_X1 U6840 ( .A1(n5943), .A2(n6475), .ZN(n5785) );
  NAND2_X1 U6841 ( .A1(n5785), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U6842 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5787) );
  MUX2_X1 U6843 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n5787), .S(n6480), .Z(n5939)
         );
  INV_X1 U6844 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9468) );
  INV_X1 U6845 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U6846 ( .A1(n5788), .A2(n5789), .ZN(n5790) );
  NAND2_X1 U6847 ( .A1(n5790), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5852) );
  XNOR2_X1 U6848 ( .A(n5852), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6269) );
  XNOR2_X1 U6849 ( .A(n5788), .B(P2_IR_REG_14__SCAN_IN), .ZN(n6257) );
  INV_X1 U6850 ( .A(n6257), .ZN(n9449) );
  NAND2_X1 U6851 ( .A1(n5791), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5795) );
  INV_X1 U6852 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U6853 ( .A1(n5795), .A2(n5792), .ZN(n5793) );
  NAND2_X1 U6854 ( .A1(n5793), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5794) );
  XNOR2_X1 U6855 ( .A(n5794), .B(P2_IR_REG_12__SCAN_IN), .ZN(n9421) );
  INV_X1 U6856 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5842) );
  OR2_X1 U6857 ( .A1(n9421), .A2(n5842), .ZN(n5844) );
  XNOR2_X1 U6858 ( .A(n5795), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8505) );
  OR2_X1 U6859 ( .A1(n5796), .A2(n5806), .ZN(n5797) );
  XNOR2_X1 U6860 ( .A(n5797), .B(n5228), .ZN(n7404) );
  OR2_X1 U6861 ( .A1(n5798), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U6862 ( .A1(n5799), .A2(n5803), .ZN(n5800) );
  OAI21_X1 U6863 ( .B1(n5802), .B2(n5800), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5801) );
  XNOR2_X1 U6864 ( .A(n5801), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U6865 ( .A1(n5802), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5825) );
  NAND2_X1 U6866 ( .A1(n5825), .A2(n5803), .ZN(n5804) );
  NAND2_X1 U6867 ( .A1(n5804), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5831) );
  NAND2_X1 U6868 ( .A1(n5798), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5805) );
  OR2_X1 U6869 ( .A1(n5807), .A2(n5806), .ZN(n5808) );
  XNOR2_X2 U6870 ( .A(n5808), .B(P2_IR_REG_4__SCAN_IN), .ZN(n10686) );
  NAND2_X1 U6871 ( .A1(n5816), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5809) );
  XNOR2_X1 U6872 ( .A(n5809), .B(P2_IR_REG_3__SCAN_IN), .ZN(n5911) );
  INV_X1 U6873 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7422) );
  OAI21_X1 U6874 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n7422), .A(n5868), .ZN(n5811) );
  NAND2_X1 U6875 ( .A1(n5871), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U6876 ( .A1(n5811), .A2(n5810), .ZN(n10663) );
  INV_X1 U6877 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10662) );
  NOR2_X1 U6878 ( .A1(n10663), .A2(n10662), .ZN(n5812) );
  AOI21_X1 U6879 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n5871), .A(n5812), .ZN(
        n7443) );
  NAND2_X1 U6880 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5813), .ZN(n5815) );
  INV_X1 U6881 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5818) );
  AOI22_X1 U6882 ( .A1(n7450), .A2(P2_REG2_REG_2__SCAN_IN), .B1(n5818), .B2(
        n7363), .ZN(n7442) );
  NOR2_X1 U6883 ( .A1(n5911), .A2(n5820), .ZN(n5821) );
  INV_X1 U6884 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n8400) );
  INV_X1 U6885 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5822) );
  AOI22_X1 U6886 ( .A1(n10686), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n5822), .B2(
        n7369), .ZN(n10679) );
  NOR2_X1 U6887 ( .A1(n10702), .A2(n5823), .ZN(n5824) );
  INV_X1 U6888 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10698) );
  INV_X1 U6889 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5826) );
  MUX2_X1 U6890 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n5826), .S(n7467), .Z(n7462)
         );
  INV_X1 U6891 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10876) );
  INV_X1 U6892 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U6893 ( .A1(n5831), .A2(n5830), .ZN(n5832) );
  NAND2_X1 U6894 ( .A1(n5832), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5834) );
  INV_X1 U6895 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U6896 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7392), .ZN(n5835) );
  OAI21_X1 U6897 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7392), .A(n5835), .ZN(
        n7846) );
  NOR2_X1 U6898 ( .A1(n6195), .A2(n5837), .ZN(n5838) );
  INV_X1 U6899 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8127) );
  XNOR2_X1 U6900 ( .A(n5837), .B(n6195), .ZN(n8128) );
  NOR2_X1 U6901 ( .A1(n8127), .A2(n8128), .ZN(n8126) );
  NAND2_X1 U6902 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7404), .ZN(n5839) );
  OAI21_X1 U6903 ( .B1(n7404), .B2(P2_REG2_REG_10__SCAN_IN), .A(n5839), .ZN(
        n8207) );
  NOR2_X1 U6904 ( .A1(n8505), .A2(n5840), .ZN(n5841) );
  INV_X1 U6905 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8499) );
  NOR2_X1 U6906 ( .A1(n5841), .A2(n8498), .ZN(n9408) );
  MUX2_X1 U6907 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n5842), .S(n9421), .Z(n9407)
         );
  NOR2_X1 U6908 ( .A1(n9408), .A2(n9407), .ZN(n9406) );
  INV_X1 U6909 ( .A(n9406), .ZN(n5843) );
  NAND2_X1 U6910 ( .A1(n5844), .A2(n5843), .ZN(n5846) );
  NAND2_X1 U6911 ( .A1(n5751), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5845) );
  XNOR2_X1 U6912 ( .A(n5845), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9442) );
  INV_X1 U6913 ( .A(n9442), .ZN(n7472) );
  INV_X1 U6914 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5847) );
  MUX2_X1 U6915 ( .A(n5847), .B(P2_REG2_REG_14__SCAN_IN), .S(n6257), .Z(n5848)
         );
  INV_X1 U6916 ( .A(n5848), .ZN(n9451) );
  XNOR2_X1 U6917 ( .A(n6269), .B(n5849), .ZN(n9469) );
  NOR2_X1 U6918 ( .A1(n6269), .A2(n5849), .ZN(n5850) );
  INV_X1 U6919 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5896) );
  INV_X1 U6920 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U6921 ( .A1(n5852), .A2(n5851), .ZN(n5853) );
  NAND2_X1 U6922 ( .A1(n5853), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5855) );
  INV_X1 U6923 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U6924 ( .A1(n5855), .A2(n5854), .ZN(n5857) );
  OR2_X1 U6925 ( .A1(n5855), .A2(n5854), .ZN(n5856) );
  MUX2_X1 U6926 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n5896), .S(n9493), .Z(n9489)
         );
  INV_X1 U6927 ( .A(n9493), .ZN(n7698) );
  NAND2_X1 U6928 ( .A1(n5857), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5858) );
  XNOR2_X1 U6929 ( .A(n5858), .B(P2_IR_REG_17__SCAN_IN), .ZN(n6297) );
  INV_X1 U6930 ( .A(n6297), .ZN(n9506) );
  INV_X1 U6931 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9501) );
  XNOR2_X1 U6932 ( .A(n5861), .B(n5741), .ZN(n9527) );
  XNOR2_X1 U6933 ( .A(n9527), .B(P2_REG2_REG_18__SCAN_IN), .ZN(n9513) );
  INV_X1 U6934 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8701) );
  INV_X1 U6935 ( .A(n9527), .ZN(n9522) );
  NOR2_X1 U6936 ( .A1(n5864), .A2(P2_U3151), .ZN(n9789) );
  AND2_X1 U6937 ( .A1(n5943), .A2(n9789), .ZN(n7425) );
  NAND2_X1 U6938 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9273) );
  INV_X1 U6939 ( .A(n7721), .ZN(n5865) );
  NOR2_X1 U6940 ( .A1(n7722), .A2(n5865), .ZN(n5866) );
  NAND2_X1 U6941 ( .A1(n9505), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5867) );
  OAI211_X1 U6942 ( .C1(n5710), .C2(n10724), .A(n9273), .B(n5867), .ZN(n5950)
         );
  INV_X1 U6943 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10716) );
  INV_X1 U6944 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7480) );
  INV_X1 U6945 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7421) );
  OAI21_X1 U6946 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n7421), .A(n5868), .ZN(n5870) );
  NAND2_X1 U6947 ( .A1(n5871), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5869) );
  INV_X1 U6948 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10664) );
  INV_X1 U6949 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7641) );
  NOR2_X1 U6950 ( .A1(n5911), .A2(n5873), .ZN(n5874) );
  AOI22_X1 U6951 ( .A1(n10686), .A2(P2_REG1_REG_4__SCAN_IN), .B1(n6131), .B2(
        n7369), .ZN(n10676) );
  NOR2_X1 U6952 ( .A1(n10702), .A2(n5875), .ZN(n5876) );
  INV_X1 U6953 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10695) );
  NOR2_X1 U6954 ( .A1(n10695), .A2(n10694), .ZN(n10693) );
  INV_X1 U6955 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7925) );
  AOI22_X1 U6956 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(n7467), .B1(n7374), .B2(
        n7925), .ZN(n7455) );
  NOR2_X1 U6957 ( .A1(n7456), .A2(n7455), .ZN(n7454) );
  XNOR2_X1 U6958 ( .A(n5877), .B(n10721), .ZN(n10715) );
  NOR2_X1 U6959 ( .A1(n10721), .A2(n5877), .ZN(n5878) );
  NAND2_X1 U6960 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7392), .ZN(n5879) );
  OAI21_X1 U6961 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7392), .A(n5879), .ZN(
        n7857) );
  NOR2_X1 U6962 ( .A1(n6195), .A2(n5880), .ZN(n5881) );
  INV_X1 U6963 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8138) );
  INV_X1 U6964 ( .A(n6195), .ZN(n8135) );
  NOR2_X1 U6965 ( .A1(n8138), .A2(n8137), .ZN(n8136) );
  NAND2_X1 U6966 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7404), .ZN(n5882) );
  OAI21_X1 U6967 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7404), .A(n5882), .ZN(
        n8199) );
  INV_X1 U6968 ( .A(n5882), .ZN(n5883) );
  INV_X1 U6969 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8497) );
  NOR2_X1 U6970 ( .A1(n8505), .A2(n5884), .ZN(n5885) );
  INV_X1 U6971 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8270) );
  INV_X1 U6972 ( .A(n9421), .ZN(n7433) );
  AOI22_X1 U6973 ( .A1(n9421), .A2(P2_REG1_REG_12__SCAN_IN), .B1(n8270), .B2(
        n7433), .ZN(n9417) );
  NOR2_X1 U6974 ( .A1(n9421), .A2(n8270), .ZN(n5886) );
  NAND2_X1 U6975 ( .A1(n5888), .A2(n7472), .ZN(n5887) );
  INV_X1 U6976 ( .A(n5887), .ZN(n5889) );
  INV_X1 U6977 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9437) );
  INV_X1 U6978 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8694) );
  AOI22_X1 U6979 ( .A1(n6257), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n8694), .B2(
        n9449), .ZN(n9445) );
  AOI21_X2 U6980 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n9449), .A(n9444), .ZN(
        n5890) );
  NOR2_X1 U6981 ( .A1(n6269), .A2(n5890), .ZN(n5891) );
  INV_X1 U6982 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9462) );
  INV_X1 U6983 ( .A(n6269), .ZN(n9466) );
  XOR2_X1 U6984 ( .A(n9466), .B(n5890), .Z(n9461) );
  INV_X1 U6985 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8778) );
  AOI22_X1 U6986 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n9493), .B1(n7698), .B2(
        n8778), .ZN(n9479) );
  NOR2_X1 U6987 ( .A1(n6297), .A2(n5098), .ZN(n5892) );
  INV_X1 U6988 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9498) );
  NAND2_X1 U6989 ( .A1(n9522), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5893) );
  OAI21_X1 U6990 ( .B1(n9522), .B2(P2_REG1_REG_18__SCAN_IN), .A(n5893), .ZN(
        n9509) );
  INV_X1 U6991 ( .A(n5893), .ZN(n5894) );
  XNOR2_X1 U6992 ( .A(n6480), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n5937) );
  XNOR2_X1 U6993 ( .A(n5895), .B(n5937), .ZN(n5948) );
  MUX2_X1 U6994 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n5088), .Z(n5933) );
  XNOR2_X1 U6995 ( .A(n5933), .B(n6297), .ZN(n9500) );
  MUX2_X1 U6996 ( .A(n5896), .B(n8778), .S(n5191), .Z(n5897) );
  NAND2_X1 U6997 ( .A1(n5897), .A2(n9493), .ZN(n5932) );
  XNOR2_X1 U6998 ( .A(n5897), .B(n7698), .ZN(n9483) );
  MUX2_X1 U6999 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n5191), .Z(n5898) );
  OR2_X1 U7000 ( .A1(n5898), .A2(n9466), .ZN(n5931) );
  XNOR2_X1 U7001 ( .A(n5898), .B(n6269), .ZN(n9465) );
  MUX2_X1 U7002 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n5088), .Z(n5899) );
  OR2_X1 U7003 ( .A1(n5899), .A2(n9449), .ZN(n5930) );
  XNOR2_X1 U7004 ( .A(n5899), .B(n6257), .ZN(n9448) );
  MUX2_X1 U7005 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n5191), .Z(n5900) );
  OR2_X1 U7006 ( .A1(n5900), .A2(n7472), .ZN(n5929) );
  XNOR2_X1 U7007 ( .A(n5900), .B(n9442), .ZN(n9431) );
  MUX2_X1 U7008 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n5088), .Z(n5901) );
  OR2_X1 U7009 ( .A1(n5901), .A2(n7433), .ZN(n5928) );
  XNOR2_X1 U7010 ( .A(n5901), .B(n9421), .ZN(n9411) );
  MUX2_X1 U7011 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n5191), .Z(n5926) );
  INV_X1 U7012 ( .A(n8505), .ZN(n7420) );
  OR2_X1 U7013 ( .A1(n5926), .A2(n7420), .ZN(n5927) );
  MUX2_X1 U7014 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n5191), .Z(n5925) );
  MUX2_X1 U7015 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n5088), .Z(n5923) );
  INV_X1 U7016 ( .A(n5923), .ZN(n5902) );
  NAND2_X1 U7017 ( .A1(n5902), .A2(n6195), .ZN(n8129) );
  INV_X1 U7018 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8515) );
  INV_X1 U7019 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5903) );
  MUX2_X1 U7020 ( .A(n8515), .B(n5903), .S(n5191), .Z(n5921) );
  INV_X1 U7021 ( .A(n7392), .ZN(n7862) );
  NAND2_X1 U7022 ( .A1(n5921), .A2(n7862), .ZN(n5920) );
  INV_X1 U7023 ( .A(n5920), .ZN(n5922) );
  MUX2_X1 U7024 ( .A(n10876), .B(n10716), .S(n5088), .Z(n5918) );
  NAND2_X1 U7025 ( .A1(n5918), .A2(n10721), .ZN(n5917) );
  INV_X1 U7026 ( .A(n5917), .ZN(n5919) );
  MUX2_X1 U7027 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n5191), .Z(n5912) );
  INV_X1 U7028 ( .A(n5912), .ZN(n5913) );
  MUX2_X1 U7029 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n5088), .Z(n5906) );
  XOR2_X1 U7030 ( .A(n5868), .B(n5906), .Z(n10660) );
  MUX2_X1 U7031 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n5191), .Z(n5905) );
  INV_X1 U7032 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5904) );
  NOR2_X1 U7033 ( .A1(n5905), .A2(n5904), .ZN(n10661) );
  INV_X1 U7034 ( .A(n5906), .ZN(n5907) );
  OAI22_X1 U7035 ( .A1(n10660), .A2(n10661), .B1(n5868), .B2(n5907), .ZN(n7437) );
  MUX2_X1 U7036 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n5191), .Z(n5908) );
  XNOR2_X1 U7037 ( .A(n5908), .B(n7450), .ZN(n7436) );
  AOI22_X1 U7038 ( .A1(n7437), .A2(n7436), .B1(n5908), .B2(n7363), .ZN(n7476)
         );
  MUX2_X1 U7039 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n5191), .Z(n5909) );
  XNOR2_X1 U7040 ( .A(n5909), .B(n5911), .ZN(n7475) );
  INV_X1 U7041 ( .A(n5909), .ZN(n5910) );
  AOI22_X1 U7042 ( .A1(n7476), .A2(n7475), .B1(n5911), .B2(n5910), .ZN(n10689)
         );
  XNOR2_X1 U7043 ( .A(n5912), .B(n10686), .ZN(n10688) );
  NAND2_X1 U7044 ( .A1(n10689), .A2(n10688), .ZN(n10687) );
  OAI21_X1 U7045 ( .B1(n10686), .B2(n5913), .A(n10687), .ZN(n10706) );
  MUX2_X1 U7046 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n5191), .Z(n5914) );
  XNOR2_X1 U7047 ( .A(n5914), .B(n10702), .ZN(n10707) );
  AOI22_X1 U7048 ( .A1(n10706), .A2(n10707), .B1(n5914), .B2(n7371), .ZN(n7458) );
  MUX2_X1 U7049 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n5191), .Z(n5915) );
  XNOR2_X1 U7050 ( .A(n5915), .B(n7467), .ZN(n7457) );
  INV_X1 U7051 ( .A(n5915), .ZN(n5916) );
  AOI22_X1 U7052 ( .A1(n7458), .A2(n7457), .B1(n7467), .B2(n5916), .ZN(n10728)
         );
  OAI21_X1 U7053 ( .B1(n5918), .B2(n10721), .A(n5917), .ZN(n10727) );
  NOR2_X1 U7054 ( .A1(n10728), .A2(n10727), .ZN(n10731) );
  NOR2_X1 U7055 ( .A1(n5919), .A2(n10731), .ZN(n7849) );
  OAI21_X1 U7056 ( .B1(n5921), .B2(n7862), .A(n5920), .ZN(n7850) );
  NOR2_X1 U7057 ( .A1(n7849), .A2(n7850), .ZN(n7851) );
  NOR2_X1 U7058 ( .A1(n5922), .A2(n7851), .ZN(n8132) );
  NAND2_X1 U7059 ( .A1(n8129), .A2(n8132), .ZN(n5924) );
  NAND2_X1 U7060 ( .A1(n5923), .A2(n8135), .ZN(n8130) );
  INV_X1 U7061 ( .A(n7404), .ZN(n8212) );
  XNOR2_X1 U7062 ( .A(n5925), .B(n8212), .ZN(n8202) );
  NAND2_X1 U7063 ( .A1(n8203), .A2(n8202), .ZN(n8201) );
  OAI21_X1 U7064 ( .B1(n5925), .B2(n7404), .A(n8201), .ZN(n8508) );
  XNOR2_X1 U7065 ( .A(n5926), .B(n8505), .ZN(n8507) );
  NAND2_X1 U7066 ( .A1(n8508), .A2(n8507), .ZN(n8506) );
  NAND2_X1 U7067 ( .A1(n5927), .A2(n8506), .ZN(n9410) );
  NAND2_X1 U7068 ( .A1(n9411), .A2(n9410), .ZN(n9409) );
  NAND2_X1 U7069 ( .A1(n5928), .A2(n9409), .ZN(n9430) );
  NAND2_X1 U7070 ( .A1(n9431), .A2(n9430), .ZN(n9429) );
  NAND2_X1 U7071 ( .A1(n5929), .A2(n9429), .ZN(n9447) );
  NAND2_X1 U7072 ( .A1(n9448), .A2(n9447), .ZN(n9446) );
  NAND2_X1 U7073 ( .A1(n5930), .A2(n9446), .ZN(n9464) );
  NAND2_X1 U7074 ( .A1(n9465), .A2(n9464), .ZN(n9463) );
  NAND2_X1 U7075 ( .A1(n5931), .A2(n9463), .ZN(n9482) );
  NAND2_X1 U7076 ( .A1(n9483), .A2(n9482), .ZN(n9481) );
  NAND2_X1 U7077 ( .A1(n5932), .A2(n9481), .ZN(n9499) );
  NOR2_X1 U7078 ( .A1(n5933), .A2(n9506), .ZN(n5934) );
  AOI21_X1 U7079 ( .B1(n9500), .B2(n9499), .A(n5934), .ZN(n5936) );
  MUX2_X1 U7080 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n5191), .Z(n5935) );
  NOR2_X1 U7081 ( .A1(n5936), .A2(n5935), .ZN(n9518) );
  NAND2_X1 U7082 ( .A1(n5936), .A2(n5935), .ZN(n9519) );
  OAI21_X1 U7083 ( .B1(n9518), .B2(n9527), .A(n9519), .ZN(n5941) );
  INV_X1 U7084 ( .A(n5937), .ZN(n5938) );
  MUX2_X1 U7085 ( .A(n5939), .B(n5938), .S(n5088), .Z(n5940) );
  XNOR2_X1 U7086 ( .A(n5941), .B(n5940), .ZN(n5946) );
  INV_X1 U7087 ( .A(n8783), .ZN(n5942) );
  INV_X1 U7088 ( .A(n5864), .ZN(n6467) );
  NOR2_X2 U7089 ( .A1(n10657), .A2(n6467), .ZN(n10729) );
  NOR2_X1 U7090 ( .A1(n5191), .A2(P2_U3151), .ZN(n8756) );
  NAND2_X1 U7091 ( .A1(n5943), .A2(n8756), .ZN(n5944) );
  MUX2_X1 U7092 ( .A(n5944), .B(n10657), .S(n6467), .Z(n9521) );
  NOR2_X1 U7093 ( .A1(n9521), .A2(n8042), .ZN(n5945) );
  NAND2_X1 U7094 ( .A1(n7312), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5964) );
  INV_X1 U7095 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9698) );
  OR2_X1 U7096 ( .A1(n5085), .A2(n9698), .ZN(n5963) );
  INV_X1 U7097 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8766) );
  NAND2_X1 U7098 ( .A1(n6141), .A2(n9116), .ZN(n6154) );
  INV_X1 U7099 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9515) );
  NAND2_X1 U7100 ( .A1(n6311), .A2(n9515), .ZN(n6324) );
  INV_X1 U7101 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9289) );
  INV_X1 U7102 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9349) );
  INV_X1 U7103 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9327) );
  INV_X1 U7104 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9296) );
  INV_X1 U7105 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9375) );
  OR2_X1 U7106 ( .A1(n6388), .A2(n9375), .ZN(n5960) );
  OR2_X1 U7107 ( .A1(n6102), .A2(n9577), .ZN(n5962) );
  INV_X1 U7108 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9754) );
  OR2_X1 U7109 ( .A1(n6470), .A2(n9754), .ZN(n5961) );
  AND2_X1 U7110 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U7111 ( .A1(n7361), .A2(n5966), .ZN(n6657) );
  AND2_X1 U7112 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U7113 ( .A1(n5974), .A2(n5967), .ZN(n6096) );
  NAND2_X1 U7114 ( .A1(n5968), .A2(SI_1_), .ZN(n5969) );
  MUX2_X1 U7115 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n5974), .Z(n5971) );
  INV_X1 U7116 ( .A(SI_2_), .ZN(n5970) );
  XNOR2_X1 U7117 ( .A(n5971), .B(n5970), .ZN(n6108) );
  NAND2_X1 U7118 ( .A1(n6107), .A2(n6108), .ZN(n5973) );
  NAND2_X1 U7119 ( .A1(n5971), .A2(SI_2_), .ZN(n5972) );
  NAND2_X1 U7120 ( .A1(n5973), .A2(n5972), .ZN(n6122) );
  MUX2_X1 U7121 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n5974), .Z(n5975) );
  INV_X1 U7122 ( .A(SI_3_), .ZN(n8883) );
  XNOR2_X1 U7123 ( .A(n5975), .B(n8883), .ZN(n6123) );
  NAND2_X1 U7124 ( .A1(n5975), .A2(SI_3_), .ZN(n5976) );
  INV_X1 U7125 ( .A(SI_4_), .ZN(n8884) );
  INV_X1 U7126 ( .A(SI_5_), .ZN(n9083) );
  NAND2_X1 U7127 ( .A1(n5979), .A2(SI_5_), .ZN(n5980) );
  MUX2_X1 U7128 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n7362), .Z(n5981) );
  INV_X1 U7129 ( .A(SI_6_), .ZN(n8878) );
  XNOR2_X1 U7130 ( .A(n5981), .B(n8878), .ZN(n6161) );
  NAND2_X1 U7131 ( .A1(n6160), .A2(n6161), .ZN(n5983) );
  NAND2_X1 U7132 ( .A1(n5981), .A2(SI_6_), .ZN(n5982) );
  MUX2_X1 U7133 ( .A(n7396), .B(n7393), .S(n7362), .Z(n5986) );
  INV_X1 U7134 ( .A(SI_8_), .ZN(n8877) );
  NAND2_X1 U7135 ( .A1(n5986), .A2(n8877), .ZN(n5989) );
  INV_X1 U7136 ( .A(n5986), .ZN(n5987) );
  NAND2_X1 U7137 ( .A1(n5987), .A2(SI_8_), .ZN(n5988) );
  NAND2_X1 U7138 ( .A1(n5989), .A2(n5988), .ZN(n6177) );
  MUX2_X1 U7139 ( .A(n9180), .B(n7399), .S(n7362), .Z(n5990) );
  NAND2_X1 U7140 ( .A1(n5990), .A2(n9077), .ZN(n5993) );
  INV_X1 U7141 ( .A(n5990), .ZN(n5991) );
  NAND2_X1 U7142 ( .A1(n5991), .A2(SI_9_), .ZN(n5992) );
  NAND2_X1 U7143 ( .A1(n6194), .A2(n5727), .ZN(n5994) );
  MUX2_X1 U7144 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n7362), .Z(n5996) );
  XNOR2_X1 U7145 ( .A(n5996), .B(n9078), .ZN(n6208) );
  INV_X1 U7146 ( .A(n6208), .ZN(n5995) );
  NAND2_X1 U7147 ( .A1(n5996), .A2(SI_10_), .ZN(n5997) );
  INV_X1 U7148 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5998) );
  MUX2_X1 U7149 ( .A(n7418), .B(n5998), .S(n7362), .Z(n6000) );
  INV_X1 U7150 ( .A(SI_11_), .ZN(n5999) );
  INV_X1 U7151 ( .A(n6000), .ZN(n6001) );
  NAND2_X1 U7152 ( .A1(n6001), .A2(SI_11_), .ZN(n6002) );
  NAND2_X1 U7153 ( .A1(n6003), .A2(n6002), .ZN(n6220) );
  MUX2_X1 U7154 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n7362), .Z(n6004) );
  MUX2_X1 U7155 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n7362), .Z(n6005) );
  XNOR2_X1 U7156 ( .A(n6005), .B(SI_13_), .ZN(n6244) );
  NAND2_X1 U7157 ( .A1(n6005), .A2(SI_13_), .ZN(n6006) );
  NAND2_X1 U7158 ( .A1(n6007), .A2(n6006), .ZN(n6256) );
  MUX2_X1 U7159 ( .A(n7559), .B(n7557), .S(n7362), .Z(n6008) );
  INV_X1 U7160 ( .A(n6008), .ZN(n6009) );
  NAND2_X1 U7161 ( .A1(n6009), .A2(SI_14_), .ZN(n6010) );
  NAND2_X1 U7162 ( .A1(n6011), .A2(n6010), .ZN(n6255) );
  MUX2_X1 U7163 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n7362), .Z(n6013) );
  INV_X1 U7164 ( .A(SI_15_), .ZN(n6012) );
  NAND2_X1 U7165 ( .A1(n6013), .A2(SI_15_), .ZN(n6014) );
  MUX2_X1 U7166 ( .A(n9169), .B(n7700), .S(n7362), .Z(n6017) );
  INV_X1 U7167 ( .A(SI_16_), .ZN(n6016) );
  INV_X1 U7168 ( .A(n6017), .ZN(n6018) );
  NAND2_X1 U7169 ( .A1(n6018), .A2(SI_16_), .ZN(n6019) );
  NAND2_X1 U7170 ( .A1(n6020), .A2(n6019), .ZN(n6282) );
  NAND2_X1 U7171 ( .A1(n6021), .A2(n6020), .ZN(n6296) );
  MUX2_X1 U7172 ( .A(n9168), .B(n7819), .S(n7362), .Z(n6022) );
  NAND2_X1 U7173 ( .A1(n6022), .A2(n9064), .ZN(n6025) );
  INV_X1 U7174 ( .A(n6022), .ZN(n6023) );
  NAND2_X1 U7175 ( .A1(n6023), .A2(SI_17_), .ZN(n6024) );
  NAND2_X1 U7176 ( .A1(n6296), .A2(n6295), .ZN(n6026) );
  MUX2_X1 U7177 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n7362), .Z(n6028) );
  INV_X1 U7178 ( .A(SI_18_), .ZN(n6027) );
  XNOR2_X1 U7179 ( .A(n6028), .B(n6027), .ZN(n6307) );
  INV_X1 U7180 ( .A(n6307), .ZN(n6030) );
  NAND2_X1 U7181 ( .A1(n6028), .A2(SI_18_), .ZN(n6029) );
  MUX2_X1 U7182 ( .A(n8041), .B(n8044), .S(n7362), .Z(n6032) );
  INV_X1 U7183 ( .A(SI_19_), .ZN(n6031) );
  NAND2_X1 U7184 ( .A1(n6032), .A2(n6031), .ZN(n6035) );
  INV_X1 U7185 ( .A(n6032), .ZN(n6033) );
  NAND2_X1 U7186 ( .A1(n6033), .A2(SI_19_), .ZN(n6034) );
  NAND2_X1 U7187 ( .A1(n6035), .A2(n6034), .ZN(n6318) );
  MUX2_X1 U7188 ( .A(n8084), .B(n8108), .S(n7362), .Z(n6036) );
  INV_X1 U7189 ( .A(SI_20_), .ZN(n9060) );
  NAND2_X1 U7190 ( .A1(n6036), .A2(n9060), .ZN(n6039) );
  INV_X1 U7191 ( .A(n6036), .ZN(n6037) );
  NAND2_X1 U7192 ( .A1(n6037), .A2(SI_20_), .ZN(n6038) );
  NAND2_X1 U7193 ( .A1(n6335), .A2(n6039), .ZN(n6345) );
  MUX2_X1 U7194 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n7362), .Z(n6040) );
  XNOR2_X1 U7195 ( .A(n6040), .B(n9059), .ZN(n6344) );
  INV_X1 U7196 ( .A(n6344), .ZN(n6042) );
  NAND2_X1 U7197 ( .A1(n6040), .A2(SI_21_), .ZN(n6041) );
  OAI21_X1 U7198 ( .B1(n6345), .B2(n6042), .A(n6041), .ZN(n6358) );
  MUX2_X1 U7199 ( .A(n9156), .B(n8264), .S(n7362), .Z(n6043) );
  INV_X1 U7200 ( .A(SI_22_), .ZN(n9055) );
  NAND2_X1 U7201 ( .A1(n6043), .A2(n9055), .ZN(n6046) );
  INV_X1 U7202 ( .A(n6043), .ZN(n6044) );
  NAND2_X1 U7203 ( .A1(n6044), .A2(SI_22_), .ZN(n6045) );
  NAND2_X1 U7204 ( .A1(n6046), .A2(n6045), .ZN(n6357) );
  MUX2_X1 U7205 ( .A(n9155), .B(n8417), .S(n7362), .Z(n6047) );
  INV_X1 U7206 ( .A(SI_23_), .ZN(n9054) );
  NAND2_X1 U7207 ( .A1(n6047), .A2(n9054), .ZN(n6051) );
  INV_X1 U7208 ( .A(n6047), .ZN(n6048) );
  NAND2_X1 U7209 ( .A1(n6048), .A2(SI_23_), .ZN(n6049) );
  NAND2_X1 U7210 ( .A1(n6051), .A2(n6049), .ZN(n6065) );
  INV_X1 U7211 ( .A(n6065), .ZN(n6050) );
  INV_X1 U7212 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8676) );
  MUX2_X1 U7213 ( .A(n9154), .B(n8676), .S(n7362), .Z(n6052) );
  INV_X1 U7214 ( .A(SI_24_), .ZN(n9050) );
  NAND2_X1 U7215 ( .A1(n6052), .A2(n9050), .ZN(n6055) );
  INV_X1 U7216 ( .A(n6052), .ZN(n6053) );
  NAND2_X1 U7217 ( .A1(n6053), .A2(SI_24_), .ZN(n6054) );
  MUX2_X1 U7218 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n7362), .Z(n6057) );
  INV_X1 U7219 ( .A(SI_25_), .ZN(n6056) );
  XNOR2_X1 U7220 ( .A(n6057), .B(n6056), .ZN(n6383) );
  INV_X1 U7221 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n6061) );
  MUX2_X1 U7222 ( .A(n9148), .B(n6061), .S(n7362), .Z(n6058) );
  INV_X1 U7223 ( .A(SI_26_), .ZN(n9037) );
  NAND2_X1 U7224 ( .A1(n6058), .A2(n9037), .ZN(n6397) );
  INV_X1 U7225 ( .A(n6058), .ZN(n6059) );
  NAND2_X1 U7226 ( .A1(n6059), .A2(SI_26_), .ZN(n6060) );
  NAND2_X1 U7227 ( .A1(n6397), .A2(n6060), .ZN(n6398) );
  INV_X2 U7228 ( .A(n6162), .ZN(n7308) );
  NAND2_X1 U7229 ( .A1(n8779), .A2(n7308), .ZN(n6063) );
  NAND2_X1 U7230 ( .A1(n6475), .A2(n7361), .ZN(n6085) );
  OR2_X1 U7231 ( .A1(n7301), .A2(n6061), .ZN(n6062) );
  NAND2_X1 U7232 ( .A1(n6066), .A2(n6065), .ZN(n6068) );
  NAND2_X1 U7233 ( .A1(n6068), .A2(n6067), .ZN(n8418) );
  NAND2_X1 U7234 ( .A1(n8418), .A2(n7308), .ZN(n6070) );
  OR2_X1 U7235 ( .A1(n6085), .A2(n8417), .ZN(n6069) );
  NAND2_X1 U7236 ( .A1(n7312), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6077) );
  INV_X1 U7237 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n6071) );
  OR2_X1 U7238 ( .A1(n6470), .A2(n6071), .ZN(n6076) );
  AND2_X1 U7239 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(n6363), .ZN(n6072) );
  NOR2_X1 U7240 ( .A1(n6377), .A2(n6072), .ZN(n9264) );
  OR2_X1 U7241 ( .A1(n6102), .A2(n9264), .ZN(n6075) );
  INV_X1 U7242 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n6073) );
  OR2_X1 U7243 ( .A1(n5086), .A2(n6073), .ZN(n6074) );
  INV_X1 U7244 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8244) );
  OR2_X1 U7245 ( .A1(n6102), .A2(n8244), .ZN(n6082) );
  INV_X1 U7246 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7247 ( .A1(n6115), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6079) );
  OR2_X1 U7248 ( .A1(n6085), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6086) );
  OAI211_X2 U7249 ( .C1(n5868), .C2(n6475), .A(n6087), .B(n6086), .ZN(n8245)
         );
  OR2_X2 U7250 ( .A1(n6098), .A2(n8245), .ZN(n7185) );
  NAND2_X1 U7251 ( .A1(n6098), .A2(n8245), .ZN(n7183) );
  NAND2_X1 U7252 ( .A1(n7185), .A2(n7183), .ZN(n7331) );
  NAND2_X1 U7253 ( .A1(n6115), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6089) );
  AND2_X1 U7254 ( .A1(n6089), .A2(n6088), .ZN(n6093) );
  INV_X1 U7255 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n8357) );
  OR2_X1 U7256 ( .A1(n6102), .A2(n8357), .ZN(n6092) );
  INV_X1 U7257 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6090) );
  OR2_X1 U7258 ( .A1(n6470), .A2(n6090), .ZN(n6091) );
  NAND2_X1 U7259 ( .A1(n7362), .A2(SI_0_), .ZN(n6095) );
  INV_X1 U7260 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7261 ( .A1(n6095), .A2(n6094), .ZN(n6097) );
  AND2_X1 U7262 ( .A1(n6097), .A2(n6096), .ZN(n9794) );
  MUX2_X1 U7263 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9794), .S(n6475), .Z(n8363) );
  NAND2_X1 U7264 ( .A1(n9405), .A2(n8363), .ZN(n7672) );
  NAND2_X1 U7265 ( .A1(n7331), .A2(n7672), .ZN(n6100) );
  INV_X1 U7266 ( .A(n8245), .ZN(n7733) );
  OR2_X1 U7267 ( .A1(n9404), .A2(n7733), .ZN(n6099) );
  NAND2_X1 U7268 ( .A1(n6100), .A2(n6099), .ZN(n7635) );
  NAND2_X1 U7269 ( .A1(n6115), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6106) );
  INV_X1 U7270 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6101) );
  OR2_X1 U7271 ( .A1(n6470), .A2(n6101), .ZN(n6105) );
  INV_X1 U7272 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8488) );
  OR2_X1 U7273 ( .A1(n6102), .A2(n8488), .ZN(n6103) );
  XNOR2_X1 U7274 ( .A(n6107), .B(n6108), .ZN(n7364) );
  OR2_X1 U7275 ( .A1(n6162), .A2(n7364), .ZN(n6111) );
  INV_X1 U7276 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7365) );
  OR2_X1 U7277 ( .A1(n7301), .A2(n7365), .ZN(n6110) );
  NAND2_X1 U7278 ( .A1(n6320), .A2(n7450), .ZN(n6109) );
  AND3_X2 U7279 ( .A1(n6111), .A2(n6110), .A3(n6109), .ZN(n7930) );
  NAND2_X1 U7280 ( .A1(n9403), .A2(n7930), .ZN(n7192) );
  NAND2_X2 U7281 ( .A1(n7191), .A2(n7192), .ZN(n7636) );
  NAND2_X1 U7282 ( .A1(n7635), .A2(n7636), .ZN(n6114) );
  INV_X1 U7283 ( .A(n7930), .ZN(n6112) );
  OR2_X1 U7284 ( .A1(n9403), .A2(n6112), .ZN(n6113) );
  NAND2_X1 U7285 ( .A1(n6115), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6121) );
  OR2_X1 U7286 ( .A1(n6102), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6119) );
  INV_X1 U7287 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6117) );
  OR2_X1 U7288 ( .A1(n6470), .A2(n6117), .ZN(n6118) );
  XNOR2_X1 U7289 ( .A(n6122), .B(n6123), .ZN(n7384) );
  OR2_X1 U7290 ( .A1(n6162), .A2(n7384), .ZN(n6125) );
  INV_X1 U7291 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7368) );
  OAI211_X1 U7292 ( .C1(n6475), .C2(n7491), .A(n6125), .B(n6124), .ZN(n7754)
         );
  NOR2_X1 U7293 ( .A1(n9402), .A2(n7754), .ZN(n6126) );
  NAND2_X1 U7294 ( .A1(n9402), .A2(n7754), .ZN(n6127) );
  NAND2_X1 U7295 ( .A1(n6115), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6135) );
  INV_X1 U7296 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6129) );
  OR2_X1 U7297 ( .A1(n6470), .A2(n6129), .ZN(n6134) );
  AND2_X1 U7298 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6130) );
  NOR2_X1 U7299 ( .A1(n6141), .A2(n6130), .ZN(n8311) );
  OR2_X1 U7300 ( .A1(n6102), .A2(n8311), .ZN(n6133) );
  INV_X1 U7301 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6131) );
  OR2_X1 U7302 ( .A1(n5086), .A2(n6131), .ZN(n6132) );
  NAND4_X1 U7303 ( .A1(n6135), .A2(n6134), .A3(n6133), .A4(n6132), .ZN(n9401)
         );
  XNOR2_X1 U7304 ( .A(n6136), .B(n6137), .ZN(n7378) );
  OR2_X1 U7305 ( .A1(n6162), .A2(n7378), .ZN(n6139) );
  INV_X1 U7306 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7370) );
  OR2_X1 U7307 ( .A1(n7301), .A2(n7370), .ZN(n6138) );
  OAI211_X1 U7308 ( .C1(n6475), .C2(n7369), .A(n6139), .B(n6138), .ZN(n7772)
         );
  NAND2_X1 U7309 ( .A1(n6115), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6146) );
  INV_X1 U7310 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6140) );
  OR2_X1 U7311 ( .A1(n6470), .A2(n6140), .ZN(n6145) );
  OR2_X1 U7312 ( .A1(n6141), .A2(n9116), .ZN(n6142) );
  AND2_X1 U7313 ( .A1(n6154), .A2(n6142), .ZN(n8348) );
  OR2_X1 U7314 ( .A1(n6102), .A2(n8348), .ZN(n6144) );
  OR2_X1 U7315 ( .A1(n5086), .A2(n10695), .ZN(n6143) );
  NAND4_X1 U7316 ( .A1(n6146), .A2(n6145), .A3(n6144), .A4(n6143), .ZN(n9400)
         );
  XNOR2_X1 U7317 ( .A(n6147), .B(n6148), .ZN(n7381) );
  OR2_X1 U7318 ( .A1(n6162), .A2(n7381), .ZN(n6150) );
  INV_X1 U7319 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7372) );
  OR2_X1 U7320 ( .A1(n7301), .A2(n7372), .ZN(n6149) );
  OAI211_X1 U7321 ( .C1(n6475), .C2(n7371), .A(n6150), .B(n6149), .ZN(n7779)
         );
  NOR2_X1 U7322 ( .A1(n9400), .A2(n7779), .ZN(n6151) );
  NAND2_X1 U7323 ( .A1(n9400), .A2(n7779), .ZN(n6152) );
  NAND2_X1 U7324 ( .A1(n6115), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6159) );
  INV_X1 U7325 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6153) );
  OR2_X1 U7326 ( .A1(n6470), .A2(n6153), .ZN(n6158) );
  NAND2_X1 U7327 ( .A1(n6154), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6155) );
  AND2_X1 U7328 ( .A1(n6167), .A2(n6155), .ZN(n8409) );
  OR2_X1 U7329 ( .A1(n6102), .A2(n8409), .ZN(n6157) );
  OR2_X1 U7330 ( .A1(n5085), .A2(n7925), .ZN(n6156) );
  NAND4_X1 U7331 ( .A1(n6159), .A2(n6158), .A3(n6157), .A4(n6156), .ZN(n9399)
         );
  XNOR2_X1 U7332 ( .A(n6160), .B(n6161), .ZN(n7375) );
  OR2_X1 U7333 ( .A1(n7375), .A2(n6162), .ZN(n6164) );
  INV_X1 U7334 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7376) );
  OR2_X1 U7335 ( .A1(n7301), .A2(n7376), .ZN(n6163) );
  OAI211_X1 U7336 ( .C1(n6475), .C2(n7374), .A(n6164), .B(n6163), .ZN(n7790)
         );
  AND2_X1 U7337 ( .A1(n9399), .A2(n7790), .ZN(n6165) );
  NAND2_X1 U7338 ( .A1(n7312), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6172) );
  INV_X1 U7339 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6166) );
  OR2_X1 U7340 ( .A1(n6470), .A2(n6166), .ZN(n6171) );
  AND2_X1 U7341 ( .A1(n6167), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6168) );
  NOR2_X1 U7342 ( .A1(n6182), .A2(n6168), .ZN(n7961) );
  OR2_X1 U7343 ( .A1(n6102), .A2(n7961), .ZN(n6170) );
  OR2_X1 U7344 ( .A1(n5086), .A2(n10716), .ZN(n6169) );
  NAND4_X1 U7345 ( .A1(n6172), .A2(n6171), .A3(n6170), .A4(n6169), .ZN(n9398)
         );
  NAND2_X1 U7346 ( .A1(n6704), .A2(n7308), .ZN(n6176) );
  AOI22_X1 U7347 ( .A1(n6321), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6320), .B2(
        n10721), .ZN(n6175) );
  OR2_X1 U7348 ( .A1(n9398), .A2(n7968), .ZN(n7223) );
  NAND2_X1 U7349 ( .A1(n9398), .A2(n7968), .ZN(n8443) );
  NAND2_X1 U7350 ( .A1(n7223), .A2(n8443), .ZN(n7884) );
  NAND2_X1 U7351 ( .A1(n7885), .A2(n7884), .ZN(n8446) );
  INV_X1 U7352 ( .A(n7968), .ZN(n10870) );
  OR2_X1 U7353 ( .A1(n9398), .A2(n10870), .ZN(n8445) );
  XNOR2_X1 U7354 ( .A(n6178), .B(n6177), .ZN(n7391) );
  NAND2_X1 U7355 ( .A1(n7391), .A2(n7308), .ZN(n6180) );
  AOI22_X1 U7356 ( .A1(n6321), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6320), .B2(
        n7862), .ZN(n6179) );
  INV_X1 U7357 ( .A(n8514), .ZN(n8452) );
  NAND2_X1 U7358 ( .A1(n7312), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6187) );
  INV_X1 U7359 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6181) );
  OR2_X1 U7360 ( .A1(n6470), .A2(n6181), .ZN(n6186) );
  NOR2_X1 U7361 ( .A1(n6182), .A2(n7848), .ZN(n6183) );
  OR2_X1 U7362 ( .A1(n6102), .A2(n5707), .ZN(n6185) );
  OR2_X1 U7363 ( .A1(n5085), .A2(n5903), .ZN(n6184) );
  NAND4_X1 U7364 ( .A1(n6187), .A2(n6186), .A3(n6185), .A4(n6184), .ZN(n9397)
         );
  OR2_X1 U7365 ( .A1(n8452), .A2(n9397), .ZN(n6189) );
  AND2_X1 U7366 ( .A1(n8445), .A2(n6189), .ZN(n6188) );
  INV_X1 U7367 ( .A(n6189), .ZN(n6191) );
  NAND2_X1 U7368 ( .A1(n8514), .A2(n9397), .ZN(n7209) );
  INV_X1 U7369 ( .A(n9397), .ZN(n6190) );
  NAND2_X1 U7370 ( .A1(n6190), .A2(n8452), .ZN(n7224) );
  NAND2_X1 U7371 ( .A1(n7209), .A2(n7224), .ZN(n8447) );
  OR2_X1 U7372 ( .A1(n6191), .A2(n8447), .ZN(n6192) );
  XNOR2_X1 U7373 ( .A(n6194), .B(n5727), .ZN(n7398) );
  NAND2_X1 U7374 ( .A1(n7398), .A2(n7308), .ZN(n6197) );
  AOI22_X1 U7375 ( .A1(n6321), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6320), .B2(
        n6195), .ZN(n6196) );
  NAND2_X1 U7376 ( .A1(n6197), .A2(n6196), .ZN(n8111) );
  NAND2_X1 U7377 ( .A1(n7312), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6204) );
  INV_X1 U7378 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n6198) );
  OR2_X1 U7379 ( .A1(n6470), .A2(n6198), .ZN(n6203) );
  OR2_X1 U7380 ( .A1(n6199), .A2(n8114), .ZN(n6200) );
  AND2_X1 U7381 ( .A1(n6212), .A2(n6200), .ZN(n8481) );
  OR2_X1 U7382 ( .A1(n6102), .A2(n8481), .ZN(n6202) );
  OR2_X1 U7383 ( .A1(n5086), .A2(n8138), .ZN(n6201) );
  NAND2_X1 U7384 ( .A1(n8111), .A2(n8449), .ZN(n7225) );
  NAND2_X1 U7385 ( .A1(n8111), .A2(n8252), .ZN(n6206) );
  XNOR2_X1 U7386 ( .A(n6207), .B(n6208), .ZN(n7400) );
  NAND2_X1 U7387 ( .A1(n7400), .A2(n7308), .ZN(n6210) );
  AOI22_X1 U7388 ( .A1(n6321), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6320), .B2(
        n8212), .ZN(n6209) );
  NAND2_X1 U7389 ( .A1(n6210), .A2(n6209), .ZN(n8290) );
  NAND2_X1 U7390 ( .A1(n7312), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6218) );
  INV_X1 U7391 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n6211) );
  OR2_X1 U7392 ( .A1(n6470), .A2(n6211), .ZN(n6217) );
  NAND2_X1 U7393 ( .A1(n6212), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6213) );
  AND2_X1 U7394 ( .A1(n6225), .A2(n6213), .ZN(n8287) );
  OR2_X1 U7395 ( .A1(n6102), .A2(n8287), .ZN(n6216) );
  INV_X1 U7396 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6214) );
  OR2_X1 U7397 ( .A1(n5086), .A2(n6214), .ZN(n6215) );
  OR2_X1 U7398 ( .A1(n8290), .A2(n8325), .ZN(n8318) );
  NAND2_X1 U7399 ( .A1(n8290), .A2(n8325), .ZN(n8320) );
  INV_X1 U7400 ( .A(n8325), .ZN(n9396) );
  OR2_X1 U7401 ( .A1(n8290), .A2(n9396), .ZN(n6219) );
  XNOR2_X1 U7402 ( .A(n6221), .B(n6220), .ZN(n7416) );
  NAND2_X1 U7403 ( .A1(n7416), .A2(n7308), .ZN(n6223) );
  AOI22_X1 U7404 ( .A1(n6321), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6320), .B2(
        n8505), .ZN(n6222) );
  NAND2_X1 U7405 ( .A1(n6223), .A2(n6222), .ZN(n8544) );
  NAND2_X1 U7406 ( .A1(n7312), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6230) );
  INV_X1 U7407 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n6224) );
  OR2_X1 U7408 ( .A1(n6470), .A2(n6224), .ZN(n6229) );
  NAND2_X1 U7409 ( .A1(n6225), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6226) );
  AND2_X1 U7410 ( .A1(n6236), .A2(n6226), .ZN(n8542) );
  OR2_X1 U7411 ( .A1(n6102), .A2(n8542), .ZN(n6228) );
  OR2_X1 U7412 ( .A1(n5086), .A2(n8497), .ZN(n6227) );
  NAND4_X1 U7413 ( .A1(n6230), .A2(n6229), .A3(n6228), .A4(n6227), .ZN(n9395)
         );
  NOR2_X1 U7414 ( .A1(n8544), .A2(n9395), .ZN(n7337) );
  NAND2_X1 U7415 ( .A1(n8544), .A2(n9395), .ZN(n7335) );
  XNOR2_X1 U7416 ( .A(n6232), .B(n6231), .ZN(n7430) );
  NAND2_X1 U7417 ( .A1(n7430), .A2(n7308), .ZN(n6234) );
  AOI22_X1 U7418 ( .A1(n6321), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6320), .B2(
        n9421), .ZN(n6233) );
  NAND2_X1 U7419 ( .A1(n7312), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6241) );
  INV_X1 U7420 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n6235) );
  OR2_X1 U7421 ( .A1(n6470), .A2(n6235), .ZN(n6240) );
  AND2_X1 U7422 ( .A1(n6236), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6237) );
  NOR2_X1 U7423 ( .A1(n6249), .A2(n6237), .ZN(n8522) );
  OR2_X1 U7424 ( .A1(n6102), .A2(n8522), .ZN(n6239) );
  OR2_X1 U7425 ( .A1(n5086), .A2(n8270), .ZN(n6238) );
  NAND4_X1 U7426 ( .A1(n6241), .A2(n6240), .A3(n6239), .A4(n6238), .ZN(n9394)
         );
  NAND2_X1 U7427 ( .A1(n8471), .A2(n9394), .ZN(n7241) );
  NAND2_X1 U7428 ( .A1(n8524), .A2(n8660), .ZN(n7240) );
  NAND2_X1 U7429 ( .A1(n7241), .A2(n7240), .ZN(n8266) );
  NAND2_X1 U7430 ( .A1(n8524), .A2(n9394), .ZN(n6242) );
  NAND2_X1 U7431 ( .A1(n6243), .A2(n6242), .ZN(n8458) );
  XNOR2_X1 U7432 ( .A(n6245), .B(n6244), .ZN(n7471) );
  NAND2_X1 U7433 ( .A1(n7471), .A2(n7308), .ZN(n6247) );
  AOI22_X1 U7434 ( .A1(n6321), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6320), .B2(
        n9442), .ZN(n6246) );
  NAND2_X1 U7435 ( .A1(n6247), .A2(n6246), .ZN(n8658) );
  NAND2_X1 U7436 ( .A1(n7312), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6254) );
  INV_X1 U7437 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n6248) );
  OR2_X1 U7438 ( .A1(n6470), .A2(n6248), .ZN(n6253) );
  OR2_X1 U7439 ( .A1(n6249), .A2(n8669), .ZN(n6250) );
  AND2_X1 U7440 ( .A1(n6250), .A2(n6261), .ZN(n8668) );
  OR2_X1 U7441 ( .A1(n6102), .A2(n8668), .ZN(n6252) );
  OR2_X1 U7442 ( .A1(n5085), .A2(n9437), .ZN(n6251) );
  OR2_X1 U7443 ( .A1(n8658), .A2(n8713), .ZN(n7176) );
  NAND2_X1 U7444 ( .A1(n8658), .A2(n8713), .ZN(n8528) );
  XNOR2_X1 U7445 ( .A(n6256), .B(n6255), .ZN(n7556) );
  NAND2_X1 U7446 ( .A1(n7556), .A2(n7308), .ZN(n6259) );
  AOI22_X1 U7447 ( .A1(n6321), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6320), .B2(
        n6257), .ZN(n6258) );
  NAND2_X1 U7448 ( .A1(n7312), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6265) );
  INV_X1 U7449 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n6260) );
  OR2_X1 U7450 ( .A1(n6470), .A2(n6260), .ZN(n6264) );
  AOI21_X1 U7451 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(n6261), .A(n6273), .ZN(
        n8714) );
  OR2_X1 U7452 ( .A1(n6102), .A2(n8714), .ZN(n6263) );
  OR2_X1 U7453 ( .A1(n5085), .A2(n8694), .ZN(n6262) );
  OR2_X1 U7454 ( .A1(n8706), .A2(n8767), .ZN(n7174) );
  NAND2_X1 U7455 ( .A1(n8706), .A2(n8767), .ZN(n6455) );
  NAND2_X1 U7456 ( .A1(n7174), .A2(n6455), .ZN(n8534) );
  INV_X1 U7457 ( .A(n8713), .ZN(n9393) );
  OR2_X1 U7458 ( .A1(n8658), .A2(n9393), .ZN(n8532) );
  AND2_X1 U7459 ( .A1(n8534), .A2(n8532), .ZN(n6266) );
  INV_X1 U7460 ( .A(n8767), .ZN(n9392) );
  XNOR2_X1 U7461 ( .A(n6268), .B(n6267), .ZN(n7642) );
  NAND2_X1 U7462 ( .A1(n7642), .A2(n7308), .ZN(n6271) );
  AOI22_X1 U7463 ( .A1(n6321), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6320), .B2(
        n6269), .ZN(n6270) );
  NAND2_X1 U7464 ( .A1(n7312), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6279) );
  INV_X1 U7465 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n6272) );
  OR2_X1 U7466 ( .A1(n6470), .A2(n6272), .ZN(n6278) );
  INV_X1 U7467 ( .A(n6273), .ZN(n6275) );
  INV_X1 U7468 ( .A(n6288), .ZN(n6274) );
  AOI21_X1 U7469 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(n6275), .A(n6274), .ZN(
        n8768) );
  OR2_X1 U7470 ( .A1(n6102), .A2(n8768), .ZN(n6277) );
  OR2_X1 U7471 ( .A1(n5085), .A2(n9462), .ZN(n6276) );
  NAND2_X1 U7472 ( .A1(n8760), .A2(n9307), .ZN(n7249) );
  NAND2_X1 U7473 ( .A1(n7175), .A2(n7249), .ZN(n8626) );
  INV_X1 U7474 ( .A(n9307), .ZN(n9391) );
  NAND2_X1 U7475 ( .A1(n8760), .A2(n9391), .ZN(n6280) );
  NAND2_X1 U7476 ( .A1(n6281), .A2(n6280), .ZN(n8680) );
  XNOR2_X1 U7477 ( .A(n6283), .B(n6282), .ZN(n7689) );
  NAND2_X1 U7478 ( .A1(n7689), .A2(n7308), .ZN(n6285) );
  AOI22_X1 U7479 ( .A1(n6321), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6320), .B2(
        n9493), .ZN(n6284) );
  NAND2_X1 U7480 ( .A1(n7312), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6292) );
  INV_X1 U7481 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n6286) );
  OR2_X1 U7482 ( .A1(n6470), .A2(n6286), .ZN(n6291) );
  AOI21_X1 U7483 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(n6288), .A(n6287), .ZN(
        n9310) );
  OR2_X1 U7484 ( .A1(n6102), .A2(n9310), .ZN(n6290) );
  OR2_X1 U7485 ( .A1(n5086), .A2(n8778), .ZN(n6289) );
  NAND2_X1 U7486 ( .A1(n9312), .A2(n8806), .ZN(n7253) );
  NAND2_X1 U7487 ( .A1(n7252), .A2(n7253), .ZN(n8681) );
  NAND2_X1 U7488 ( .A1(n8680), .A2(n8681), .ZN(n6294) );
  INV_X1 U7489 ( .A(n8806), .ZN(n9390) );
  NAND2_X1 U7490 ( .A1(n9312), .A2(n9390), .ZN(n6293) );
  XNOR2_X1 U7491 ( .A(n6296), .B(n6295), .ZN(n7817) );
  NAND2_X1 U7492 ( .A1(n7817), .A2(n7308), .ZN(n6299) );
  AOI22_X1 U7493 ( .A1(n6321), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6320), .B2(
        n6297), .ZN(n6298) );
  NAND2_X1 U7494 ( .A1(n7312), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6306) );
  INV_X1 U7495 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n6300) );
  OR2_X1 U7496 ( .A1(n6470), .A2(n6300), .ZN(n6305) );
  AND2_X1 U7497 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(n6301), .ZN(n6302) );
  NOR2_X1 U7498 ( .A1(n6311), .A2(n6302), .ZN(n9319) );
  OR2_X1 U7499 ( .A1(n6102), .A2(n9319), .ZN(n6304) );
  OR2_X1 U7500 ( .A1(n5086), .A2(n9498), .ZN(n6303) );
  XNOR2_X1 U7501 ( .A(n9321), .B(n8809), .ZN(n8725) );
  INV_X1 U7502 ( .A(n8809), .ZN(n9389) );
  XNOR2_X1 U7503 ( .A(n6308), .B(n6307), .ZN(n7821) );
  NAND2_X1 U7504 ( .A1(n7821), .A2(n7308), .ZN(n6310) );
  AOI22_X1 U7505 ( .A1(n6321), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6320), .B2(
        n9527), .ZN(n6309) );
  NAND2_X1 U7506 ( .A1(n7312), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6316) );
  INV_X1 U7507 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9777) );
  OR2_X1 U7508 ( .A1(n6470), .A2(n9777), .ZN(n6315) );
  OR2_X1 U7509 ( .A1(n6311), .A2(n9515), .ZN(n6312) );
  AND2_X1 U7510 ( .A1(n6312), .A2(n6324), .ZN(n9360) );
  OR2_X1 U7511 ( .A1(n6102), .A2(n9360), .ZN(n6314) );
  INV_X1 U7512 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9736) );
  OR2_X1 U7513 ( .A1(n5085), .A2(n9736), .ZN(n6313) );
  NAND4_X1 U7514 ( .A1(n6316), .A2(n6315), .A3(n6314), .A4(n6313), .ZN(n9666)
         );
  AND2_X1 U7515 ( .A1(n8811), .A2(n9666), .ZN(n6317) );
  XNOR2_X1 U7516 ( .A(n6319), .B(n6318), .ZN(n8040) );
  NAND2_X1 U7517 ( .A1(n8040), .A2(n7308), .ZN(n6323) );
  AOI22_X1 U7518 ( .A1(n6321), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6480), .B2(
        n6320), .ZN(n6322) );
  NAND2_X1 U7519 ( .A1(n7312), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6329) );
  INV_X1 U7520 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9773) );
  OR2_X1 U7521 ( .A1(n6470), .A2(n9773), .ZN(n6328) );
  NAND2_X1 U7522 ( .A1(n6324), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6325) );
  AND2_X1 U7523 ( .A1(n6338), .A2(n6325), .ZN(n9272) );
  OR2_X1 U7524 ( .A1(n6102), .A2(n9272), .ZN(n6327) );
  INV_X1 U7525 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9730) );
  OR2_X1 U7526 ( .A1(n5085), .A2(n9730), .ZN(n6326) );
  NAND2_X1 U7527 ( .A1(n9674), .A2(n9655), .ZN(n7258) );
  INV_X1 U7528 ( .A(n9655), .ZN(n9388) );
  NAND2_X1 U7529 ( .A1(n9674), .A2(n9388), .ZN(n6331) );
  OR2_X1 U7530 ( .A1(n6333), .A2(n6332), .ZN(n6334) );
  NAND2_X1 U7531 ( .A1(n6335), .A2(n6334), .ZN(n8106) );
  NAND2_X1 U7532 ( .A1(n8106), .A2(n7308), .ZN(n6337) );
  OR2_X1 U7533 ( .A1(n7301), .A2(n8108), .ZN(n6336) );
  NAND2_X1 U7534 ( .A1(n7312), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6343) );
  INV_X1 U7535 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9769) );
  OR2_X1 U7536 ( .A1(n6470), .A2(n9769), .ZN(n6342) );
  AND2_X1 U7537 ( .A1(n6338), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6339) );
  NOR2_X1 U7538 ( .A1(n6349), .A2(n6339), .ZN(n9340) );
  OR2_X1 U7539 ( .A1(n6102), .A2(n9340), .ZN(n6341) );
  INV_X1 U7540 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9726) );
  OR2_X1 U7541 ( .A1(n5086), .A2(n9726), .ZN(n6340) );
  NAND2_X1 U7542 ( .A1(n9657), .A2(n9636), .ZN(n7267) );
  INV_X1 U7543 ( .A(n9636), .ZN(n9669) );
  XNOR2_X1 U7544 ( .A(n6345), .B(n6344), .ZN(n8120) );
  NAND2_X1 U7545 ( .A1(n8120), .A2(n7308), .ZN(n6347) );
  INV_X1 U7546 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8121) );
  OR2_X1 U7547 ( .A1(n6085), .A2(n8121), .ZN(n6346) );
  NAND2_X1 U7548 ( .A1(n7312), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6356) );
  INV_X1 U7549 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n6348) );
  OR2_X1 U7550 ( .A1(n5086), .A2(n6348), .ZN(n6355) );
  NOR2_X1 U7551 ( .A1(n6349), .A2(n9289), .ZN(n6350) );
  OR2_X1 U7552 ( .A1(n6362), .A2(n6350), .ZN(n9645) );
  INV_X1 U7553 ( .A(n9645), .ZN(n6351) );
  INV_X1 U7554 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n6352) );
  OR2_X1 U7555 ( .A1(n6470), .A2(n6352), .ZN(n6353) );
  NAND2_X1 U7556 ( .A1(n9719), .A2(n9654), .ZN(n7272) );
  NAND2_X1 U7557 ( .A1(n7271), .A2(n7272), .ZN(n9634) );
  INV_X1 U7558 ( .A(n9719), .ZN(n9648) );
  XNOR2_X1 U7559 ( .A(n6358), .B(n6357), .ZN(n8261) );
  NAND2_X1 U7560 ( .A1(n8261), .A2(n7308), .ZN(n6360) );
  OR2_X1 U7561 ( .A1(n7301), .A2(n8264), .ZN(n6359) );
  NAND2_X1 U7562 ( .A1(n7312), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6369) );
  INV_X1 U7563 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n6361) );
  OR2_X1 U7564 ( .A1(n6470), .A2(n6361), .ZN(n6368) );
  OR2_X1 U7565 ( .A1(n6362), .A2(n9349), .ZN(n6364) );
  AND2_X1 U7566 ( .A1(n6364), .A2(n6363), .ZN(n9624) );
  OR2_X1 U7567 ( .A1(n6102), .A2(n9624), .ZN(n6367) );
  INV_X1 U7568 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6365) );
  OR2_X1 U7569 ( .A1(n5085), .A2(n6365), .ZN(n6366) );
  NAND2_X1 U7570 ( .A1(n8820), .A2(n9638), .ZN(n6370) );
  OAI21_X1 U7571 ( .B1(n9618), .B2(n9601), .A(n9610), .ZN(n6372) );
  XNOR2_X1 U7572 ( .A(n6374), .B(n6373), .ZN(n8586) );
  NAND2_X1 U7573 ( .A1(n8586), .A2(n7308), .ZN(n6376) );
  OR2_X1 U7574 ( .A1(n6085), .A2(n8676), .ZN(n6375) );
  NAND2_X1 U7575 ( .A1(n7312), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6382) );
  INV_X1 U7576 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9762) );
  OR2_X1 U7577 ( .A1(n6470), .A2(n9762), .ZN(n6381) );
  NOR2_X1 U7578 ( .A1(n6377), .A2(n9327), .ZN(n6378) );
  OR2_X1 U7579 ( .A1(n6386), .A2(n6378), .ZN(n9605) );
  INV_X1 U7580 ( .A(n9605), .ZN(n9332) );
  INV_X1 U7581 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9708) );
  OR2_X1 U7582 ( .A1(n5085), .A2(n9708), .ZN(n6379) );
  INV_X1 U7583 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8633) );
  OR2_X1 U7584 ( .A1(n7301), .A2(n8633), .ZN(n6385) );
  NAND2_X1 U7585 ( .A1(n7312), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6392) );
  INV_X1 U7586 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9758) );
  OR2_X1 U7587 ( .A1(n6470), .A2(n9758), .ZN(n6391) );
  NOR2_X1 U7588 ( .A1(n6386), .A2(n9296), .ZN(n6387) );
  NOR2_X1 U7589 ( .A1(n6388), .A2(n6387), .ZN(n9591) );
  OR2_X1 U7590 ( .A1(n6102), .A2(n9591), .ZN(n6390) );
  INV_X1 U7591 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9704) );
  OR2_X1 U7592 ( .A1(n5085), .A2(n9704), .ZN(n6389) );
  INV_X1 U7593 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9149) );
  INV_X1 U7594 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6403) );
  MUX2_X1 U7595 ( .A(n9149), .B(n6403), .S(n7362), .Z(n6400) );
  INV_X1 U7596 ( .A(SI_27_), .ZN(n9039) );
  NAND2_X1 U7597 ( .A1(n6400), .A2(n9039), .ZN(n6414) );
  INV_X1 U7598 ( .A(n6400), .ZN(n6401) );
  NAND2_X1 U7599 ( .A1(n6401), .A2(SI_27_), .ZN(n6402) );
  NAND2_X1 U7600 ( .A1(n8755), .A2(n7308), .ZN(n6405) );
  OR2_X1 U7601 ( .A1(n6085), .A2(n6403), .ZN(n6404) );
  NAND2_X1 U7602 ( .A1(n7312), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6410) );
  INV_X1 U7603 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9750) );
  OR2_X1 U7604 ( .A1(n6470), .A2(n9750), .ZN(n6409) );
  XNOR2_X1 U7605 ( .A(P2_REG3_REG_27__SCAN_IN), .B(n6406), .ZN(n9568) );
  OR2_X1 U7606 ( .A1(n6102), .A2(n9568), .ZN(n6408) );
  INV_X1 U7607 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9692) );
  OR2_X1 U7608 ( .A1(n5086), .A2(n9692), .ZN(n6407) );
  NAND4_X2 U7609 ( .A1(n6410), .A2(n6409), .A3(n6408), .A4(n6407), .ZN(n9385)
         );
  NAND2_X1 U7610 ( .A1(n8841), .A2(n9385), .ZN(n6411) );
  INV_X2 U7611 ( .A(n9385), .ZN(n9576) );
  AOI21_X1 U7612 ( .B1(n9561), .B2(n6411), .A(n5723), .ZN(n9549) );
  NAND2_X1 U7613 ( .A1(n6413), .A2(n6412), .ZN(n6415) );
  MUX2_X1 U7614 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n7362), .Z(n6433) );
  INV_X1 U7615 ( .A(SI_28_), .ZN(n9038) );
  XNOR2_X1 U7616 ( .A(n6433), .B(n9038), .ZN(n6431) );
  NAND2_X1 U7617 ( .A1(n8787), .A2(n7308), .ZN(n6418) );
  INV_X1 U7618 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6416) );
  OR2_X1 U7619 ( .A1(n7301), .A2(n6416), .ZN(n6417) );
  NAND2_X1 U7620 ( .A1(n7312), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6426) );
  INV_X1 U7621 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9109) );
  NAND2_X1 U7622 ( .A1(n6420), .A2(n9109), .ZN(n9533) );
  INV_X1 U7623 ( .A(n6420), .ZN(n6421) );
  NAND2_X1 U7624 ( .A1(n6421), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6422) );
  OR2_X1 U7625 ( .A1(n6102), .A2(n9281), .ZN(n6425) );
  INV_X1 U7626 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9688) );
  OR2_X1 U7627 ( .A1(n5086), .A2(n9688), .ZN(n6424) );
  INV_X1 U7628 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9746) );
  OR2_X1 U7629 ( .A1(n6470), .A2(n9746), .ZN(n6423) );
  NAND2_X1 U7630 ( .A1(n9748), .A2(n10659), .ZN(n6427) );
  NAND2_X1 U7631 ( .A1(n9549), .A2(n6427), .ZN(n6430) );
  INV_X1 U7632 ( .A(n10659), .ZN(n6428) );
  NAND2_X1 U7633 ( .A1(n9555), .A2(n6428), .ZN(n6429) );
  NAND2_X1 U7634 ( .A1(n6430), .A2(n6429), .ZN(n6445) );
  NAND2_X1 U7635 ( .A1(n6432), .A2(n6431), .ZN(n6436) );
  INV_X1 U7636 ( .A(n6433), .ZN(n6434) );
  NAND2_X1 U7637 ( .A1(n6434), .A2(n9038), .ZN(n6435) );
  INV_X1 U7638 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8792) );
  INV_X1 U7639 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9255) );
  MUX2_X1 U7640 ( .A(n8792), .B(n9255), .S(n7362), .Z(n6547) );
  NAND2_X1 U7641 ( .A1(n8789), .A2(n7308), .ZN(n6438) );
  OR2_X1 U7642 ( .A1(n6085), .A2(n9255), .ZN(n6437) );
  INV_X1 U7643 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6439) );
  OR2_X1 U7644 ( .A1(n6128), .A2(n6439), .ZN(n6444) );
  INV_X1 U7645 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6440) );
  OR2_X1 U7646 ( .A1(n6116), .A2(n6440), .ZN(n6443) );
  INV_X1 U7647 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6441) );
  OR2_X1 U7648 ( .A1(n6470), .A2(n6441), .ZN(n6442) );
  NAND2_X1 U7649 ( .A1(n6510), .A2(n9550), .ZN(n7322) );
  XNOR2_X1 U7650 ( .A(n6445), .B(n5384), .ZN(n6479) );
  XNOR2_X1 U7651 ( .A(n6446), .B(P2_IR_REG_20__SCAN_IN), .ZN(n6465) );
  NAND2_X1 U7652 ( .A1(n7730), .A2(n6465), .ZN(n7731) );
  NAND2_X1 U7653 ( .A1(n6480), .A2(n7354), .ZN(n6504) );
  INV_X1 U7654 ( .A(n7331), .ZN(n6449) );
  INV_X1 U7655 ( .A(n8363), .ZN(n7889) );
  NAND2_X1 U7656 ( .A1(n6447), .A2(n8363), .ZN(n7736) );
  INV_X1 U7657 ( .A(n7736), .ZN(n6448) );
  NAND2_X1 U7658 ( .A1(n7671), .A2(n7185), .ZN(n7634) );
  OR2_X1 U7659 ( .A1(n9402), .A2(n8401), .ZN(n7213) );
  NAND2_X1 U7660 ( .A1(n9401), .A2(n8312), .ZN(n7179) );
  AND2_X1 U7661 ( .A1(n7200), .A2(n7179), .ZN(n7682) );
  INV_X1 U7662 ( .A(n7779), .ZN(n8349) );
  OR2_X1 U7663 ( .A1(n9400), .A2(n8349), .ZN(n7917) );
  NAND2_X1 U7664 ( .A1(n9400), .A2(n8349), .ZN(n7202) );
  INV_X1 U7665 ( .A(n7790), .ZN(n8408) );
  OR2_X1 U7666 ( .A1(n9399), .A2(n8408), .ZN(n7203) );
  NAND2_X1 U7667 ( .A1(n9399), .A2(n8408), .ZN(n7201) );
  NAND2_X1 U7668 ( .A1(n7883), .A2(n6451), .ZN(n7882) );
  AND2_X1 U7669 ( .A1(n7209), .A2(n8443), .ZN(n7219) );
  NAND2_X1 U7670 ( .A1(n8544), .A2(n8473), .ZN(n6452) );
  AND2_X1 U7671 ( .A1(n6452), .A2(n8320), .ZN(n7236) );
  NAND2_X1 U7672 ( .A1(n8100), .A2(n7236), .ZN(n6453) );
  OR2_X1 U7673 ( .A1(n8544), .A2(n8473), .ZN(n7234) );
  INV_X1 U7674 ( .A(n8266), .ZN(n6454) );
  INV_X1 U7675 ( .A(n8534), .ZN(n8529) );
  INV_X1 U7676 ( .A(n6455), .ZN(n8622) );
  NOR2_X1 U7677 ( .A1(n8626), .A2(n8622), .ZN(n6456) );
  NAND2_X1 U7678 ( .A1(n8624), .A2(n7175), .ZN(n8679) );
  INV_X1 U7679 ( .A(n8681), .ZN(n8678) );
  NAND2_X1 U7680 ( .A1(n8679), .A2(n8678), .ZN(n6457) );
  NAND2_X1 U7681 ( .A1(n6457), .A2(n7252), .ZN(n8724) );
  INV_X1 U7682 ( .A(n8725), .ZN(n6458) );
  NAND2_X1 U7683 ( .A1(n9321), .A2(n8809), .ZN(n6459) );
  NAND2_X1 U7684 ( .A1(n8811), .A2(n9316), .ZN(n7260) );
  INV_X1 U7685 ( .A(n9634), .ZN(n9641) );
  NAND2_X1 U7686 ( .A1(n9642), .A2(n9641), .ZN(n9644) );
  NAND2_X1 U7687 ( .A1(n9644), .A2(n7271), .ZN(n9628) );
  XNOR2_X1 U7688 ( .A(n9714), .B(n9611), .ZN(n9627) );
  OR2_X1 U7689 ( .A1(n9714), .A2(n9638), .ZN(n7168) );
  AND2_X1 U7690 ( .A1(n9618), .A2(n9622), .ZN(n7280) );
  NAND2_X1 U7691 ( .A1(n9710), .A2(n9601), .ZN(n7167) );
  NAND2_X1 U7692 ( .A1(n6461), .A2(n7279), .ZN(n9595) );
  NAND2_X1 U7693 ( .A1(n9702), .A2(n7285), .ZN(n9580) );
  NAND2_X1 U7694 ( .A1(n9580), .A2(n9579), .ZN(n9696) );
  OR2_X1 U7695 ( .A1(n9584), .A2(n9589), .ZN(n6462) );
  NOR2_X1 U7696 ( .A1(n8841), .A2(n9576), .ZN(n7296) );
  NAND2_X1 U7697 ( .A1(n8841), .A2(n9576), .ZN(n7292) );
  OR2_X1 U7698 ( .A1(n9555), .A2(n10659), .ZN(n6463) );
  AOI21_X1 U7699 ( .B1(n6465), .B2(n8262), .A(n6480), .ZN(n6464) );
  AND2_X1 U7700 ( .A1(n8726), .A2(n6464), .ZN(n6466) );
  NAND2_X1 U7701 ( .A1(n6481), .A2(n8042), .ZN(n6523) );
  NAND2_X1 U7702 ( .A1(n6467), .A2(n7353), .ZN(n6468) );
  NAND2_X1 U7703 ( .A1(n6475), .A2(n6468), .ZN(n7749) );
  NAND2_X1 U7704 ( .A1(n7312), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6474) );
  INV_X1 U7705 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6469) );
  OR2_X1 U7706 ( .A1(n6470), .A2(n6469), .ZN(n6473) );
  INV_X1 U7707 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6471) );
  OR2_X1 U7708 ( .A1(n5085), .A2(n6471), .ZN(n6472) );
  NAND4_X1 U7709 ( .A1(n7318), .A2(n6474), .A3(n6473), .A4(n6472), .ZN(n9384)
         );
  AND2_X1 U7710 ( .A1(n6475), .A2(P2_B_REG_SCAN_IN), .ZN(n6476) );
  NOR2_X1 U7711 ( .A1(n9637), .A2(n6476), .ZN(n9534) );
  NAND2_X1 U7712 ( .A1(n9384), .A2(n9534), .ZN(n6477) );
  OAI21_X1 U7713 ( .B1(n10659), .B2(n9635), .A(n6477), .ZN(n6478) );
  NAND2_X1 U7714 ( .A1(n6481), .A2(n6480), .ZN(n7729) );
  OR2_X1 U7715 ( .A1(n7729), .A2(n7354), .ZN(n7630) );
  XNOR2_X1 U7716 ( .A(n6484), .B(P2_B_REG_SCAN_IN), .ZN(n6486) );
  NAND2_X1 U7717 ( .A1(n6486), .A2(n6485), .ZN(n6487) );
  NAND2_X1 U7718 ( .A1(n6484), .A2(n8784), .ZN(n6489) );
  NAND2_X1 U7719 ( .A1(n6485), .A2(n8784), .ZN(n6491) );
  NAND2_X1 U7720 ( .A1(n8235), .A2(n8238), .ZN(n6520) );
  NOR2_X1 U7721 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6496) );
  NOR4_X1 U7722 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6495) );
  NOR4_X1 U7723 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6494) );
  NOR4_X1 U7724 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6493) );
  NAND4_X1 U7725 ( .A1(n6496), .A2(n6495), .A3(n6494), .A4(n6493), .ZN(n6502)
         );
  NOR4_X1 U7726 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6500) );
  NOR4_X1 U7727 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6499) );
  NOR4_X1 U7728 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6498) );
  NOR4_X1 U7729 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6497) );
  NAND4_X1 U7730 ( .A1(n6500), .A2(n6499), .A3(n6498), .A4(n6497), .ZN(n6501)
         );
  NOR2_X1 U7731 ( .A1(n6502), .A2(n6501), .ZN(n6503) );
  OR2_X1 U7732 ( .A1(n6490), .A2(n6503), .ZN(n6518) );
  OR2_X1 U7733 ( .A1(n6520), .A2(n6505), .ZN(n7746) );
  OR3_X1 U7734 ( .A1(n7730), .A2(n6481), .A3(n6504), .ZN(n7719) );
  AND2_X1 U7735 ( .A1(n8355), .A2(n7719), .ZN(n6509) );
  NOR2_X1 U7736 ( .A1(n8238), .A2(n6505), .ZN(n6506) );
  INV_X1 U7737 ( .A(n8235), .ZN(n6522) );
  NAND2_X1 U7738 ( .A1(n6506), .A2(n6522), .ZN(n7748) );
  NAND3_X1 U7739 ( .A1(n7306), .A2(n8726), .A3(n7719), .ZN(n6507) );
  INV_X1 U7740 ( .A(n7729), .ZN(n8243) );
  OR2_X1 U7741 ( .A1(n8726), .A2(n8243), .ZN(n9592) );
  AND2_X1 U7742 ( .A1(n6507), .A2(n9592), .ZN(n7717) );
  OR2_X1 U7743 ( .A1(n7748), .A2(n7717), .ZN(n6508) );
  NAND2_X1 U7744 ( .A1(n6517), .A2(n11017), .ZN(n6516) );
  NAND2_X1 U7745 ( .A1(n7397), .A2(n9720), .ZN(n7745) );
  INV_X1 U7746 ( .A(n7745), .ZN(n6511) );
  OR2_X1 U7747 ( .A1(n11017), .A2(n6441), .ZN(n6513) );
  OAI21_X1 U7748 ( .B1(n9542), .B2(n9779), .A(n6513), .ZN(n6514) );
  INV_X1 U7749 ( .A(n6514), .ZN(n6515) );
  AND2_X1 U7750 ( .A1(n6518), .A2(n7397), .ZN(n6519) );
  NOR2_X1 U7751 ( .A1(n7630), .A2(n7730), .ZN(n6521) );
  OR2_X1 U7752 ( .A1(n6522), .A2(n6521), .ZN(n6527) );
  INV_X1 U7753 ( .A(n6523), .ZN(n6524) );
  NAND3_X1 U7754 ( .A1(n6465), .A2(n7354), .A3(n8042), .ZN(n6525) );
  NAND2_X1 U7755 ( .A1(n7306), .A2(n6525), .ZN(n8236) );
  NAND2_X1 U7756 ( .A1(n7725), .A2(n8236), .ZN(n8233) );
  INV_X1 U7757 ( .A(n8238), .ZN(n6526) );
  AOI22_X1 U7758 ( .A1(n6527), .A2(n8233), .B1(n6526), .B2(n8236), .ZN(n6528)
         );
  INV_X1 U7759 ( .A(n6510), .ZN(n9542) );
  NAND2_X1 U7760 ( .A1(n6532), .A2(n6531), .ZN(P2_U3488) );
  INV_X1 U7761 ( .A(n6687), .ZN(n6534) );
  NAND2_X1 U7762 ( .A1(n6534), .A2(n6533), .ZN(n6689) );
  NAND2_X1 U7763 ( .A1(n6850), .A2(n9212), .ZN(n6537) );
  OAI21_X1 U7764 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6538) );
  NAND2_X1 U7765 ( .A1(n6987), .A2(n9221), .ZN(n6545) );
  NAND2_X1 U7766 ( .A1(n6546), .A2(n9009), .ZN(n7146) );
  NAND2_X2 U7767 ( .A1(n7950), .A2(n5452), .ZN(n7547) );
  INV_X1 U7768 ( .A(SI_29_), .ZN(n9044) );
  INV_X1 U7769 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10585) );
  INV_X1 U7770 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9260) );
  MUX2_X1 U7771 ( .A(n10585), .B(n9260), .S(n7362), .Z(n6550) );
  INV_X1 U7772 ( .A(SI_30_), .ZN(n8843) );
  NAND2_X1 U7773 ( .A1(n6550), .A2(n8843), .ZN(n6977) );
  INV_X1 U7774 ( .A(n6550), .ZN(n6551) );
  NAND2_X1 U7775 ( .A1(n6551), .A2(SI_30_), .ZN(n6552) );
  NAND2_X1 U7776 ( .A1(n6977), .A2(n6552), .ZN(n6978) );
  NAND2_X1 U7777 ( .A1(n9258), .A2(n6890), .ZN(n6558) );
  OR2_X1 U7778 ( .A1(n5092), .A2(n10585), .ZN(n6557) );
  XNOR2_X2 U7779 ( .A(n6561), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6574) );
  NAND2_X1 U7780 ( .A1(n6562), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U7781 ( .A1(n6853), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6567) );
  INV_X1 U7782 ( .A(n6668), .ZN(n6682) );
  NAND2_X1 U7783 ( .A1(n6794), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6566) );
  INV_X1 U7784 ( .A(n6574), .ZN(n10584) );
  NAND2_X1 U7785 ( .A1(n6898), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6565) );
  AND3_X1 U7786 ( .A1(n6567), .A2(n6566), .A3(n6565), .ZN(n10250) );
  NOR2_X1 U7787 ( .A1(n10226), .A2(n10250), .ZN(n7038) );
  INV_X1 U7788 ( .A(n7038), .ZN(n7129) );
  NAND2_X1 U7789 ( .A1(n6853), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6570) );
  NAND2_X1 U7790 ( .A1(n6794), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6569) );
  NAND2_X1 U7791 ( .A1(n6898), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6568) );
  NAND3_X1 U7792 ( .A1(n6570), .A2(n6569), .A3(n6568), .ZN(n10091) );
  INV_X1 U7793 ( .A(n10091), .ZN(n10230) );
  OR2_X1 U7794 ( .A1(n7129), .A2(n10230), .ZN(n7036) );
  NAND2_X1 U7795 ( .A1(n8789), .A2(n6890), .ZN(n6572) );
  OR2_X1 U7796 ( .A1(n6692), .A2(n8792), .ZN(n6571) );
  NAND2_X1 U7797 ( .A1(n6853), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6584) );
  NAND2_X1 U7798 ( .A1(n6898), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6583) );
  INV_X1 U7799 ( .A(n8790), .ZN(n6573) );
  AND2_X2 U7800 ( .A1(n6574), .A2(n6573), .ZN(n6681) );
  NAND2_X1 U7801 ( .A1(n6720), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6719) );
  NAND2_X1 U7802 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n6575) );
  NOR2_X1 U7803 ( .A1(n6719), .A2(n6575), .ZN(n6731) );
  NAND2_X1 U7804 ( .A1(n6731), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6773) );
  NAND2_X1 U7805 ( .A1(n6812), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6829) );
  INV_X1 U7806 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6828) );
  INV_X1 U7807 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6843) );
  INV_X1 U7808 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6854) );
  NAND2_X1 U7809 ( .A1(n6870), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6882) );
  INV_X1 U7810 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6881) );
  INV_X1 U7811 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6899) );
  INV_X1 U7812 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n10051) );
  NAND2_X1 U7813 ( .A1(n6627), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6601) );
  INV_X1 U7814 ( .A(n6601), .ZN(n6576) );
  NAND2_X1 U7815 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n6576), .ZN(n6927) );
  INV_X1 U7816 ( .A(n6927), .ZN(n6577) );
  NAND2_X1 U7817 ( .A1(n6577), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6942) );
  INV_X1 U7818 ( .A(n6942), .ZN(n6578) );
  NAND2_X1 U7819 ( .A1(n6578), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6953) );
  INV_X1 U7820 ( .A(n6953), .ZN(n6579) );
  NAND2_X1 U7821 ( .A1(n6579), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6955) );
  INV_X1 U7822 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6580) );
  NOR2_X1 U7823 ( .A1(n6955), .A2(n6580), .ZN(n10276) );
  NAND2_X1 U7824 ( .A1(n6956), .A2(n10276), .ZN(n6582) );
  NAND2_X1 U7825 ( .A1(n5091), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6581) );
  NAND2_X1 U7826 ( .A1(n10491), .A2(n9960), .ZN(n7125) );
  MUX2_X1 U7827 ( .A(n7125), .B(n7039), .S(n7547), .Z(n6973) );
  NAND2_X1 U7828 ( .A1(n8787), .A2(n6890), .ZN(n6586) );
  INV_X1 U7829 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10658) );
  OR2_X1 U7830 ( .A1(n5092), .A2(n10658), .ZN(n6585) );
  NAND2_X1 U7831 ( .A1(n6951), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6590) );
  NAND2_X1 U7832 ( .A1(n6898), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6589) );
  XNOR2_X1 U7833 ( .A(n6955), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n10288) );
  NAND2_X1 U7834 ( .A1(n6956), .A2(n10288), .ZN(n6588) );
  NAND2_X1 U7835 ( .A1(n5091), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6587) );
  NAND4_X1 U7836 ( .A1(n6590), .A2(n6589), .A3(n6588), .A4(n6587), .ZN(n10271)
         );
  OR2_X1 U7837 ( .A1(n10495), .A2(n10306), .ZN(n6965) );
  NAND2_X1 U7838 ( .A1(n7039), .A2(n6965), .ZN(n7127) );
  NAND2_X1 U7839 ( .A1(n7127), .A2(n6976), .ZN(n6971) );
  NAND2_X1 U7840 ( .A1(n8586), .A2(n6890), .ZN(n6592) );
  OR2_X1 U7841 ( .A1(n6692), .A2(n9154), .ZN(n6591) );
  NAND2_X2 U7842 ( .A1(n6592), .A2(n6591), .ZN(n10514) );
  NAND2_X1 U7843 ( .A1(n6951), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U7844 ( .A1(n6898), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6597) );
  INV_X1 U7845 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6593) );
  NAND2_X1 U7846 ( .A1(n6593), .A2(n6601), .ZN(n6594) );
  AND2_X1 U7847 ( .A1(n6594), .A2(n6927), .ZN(n10345) );
  NAND2_X1 U7848 ( .A1(n6956), .A2(n10345), .ZN(n6596) );
  NAND2_X1 U7849 ( .A1(n5091), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U7850 ( .A1(n10514), .A2(n9986), .ZN(n7027) );
  NAND2_X1 U7851 ( .A1(n10239), .A2(n7027), .ZN(n10342) );
  NAND2_X1 U7852 ( .A1(n8418), .A2(n6890), .ZN(n6600) );
  OR2_X1 U7853 ( .A1(n5092), .A2(n9155), .ZN(n6599) );
  NAND2_X1 U7854 ( .A1(n6898), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U7855 ( .A1(n6951), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6605) );
  OAI21_X1 U7856 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n6627), .A(n6601), .ZN(
        n6602) );
  INV_X1 U7857 ( .A(n6602), .ZN(n10358) );
  NAND2_X1 U7858 ( .A1(n6956), .A2(n10358), .ZN(n6604) );
  NAND2_X1 U7859 ( .A1(n6794), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6603) );
  NAND4_X1 U7860 ( .A1(n6606), .A2(n6605), .A3(n6604), .A4(n6603), .ZN(n10380)
         );
  INV_X1 U7861 ( .A(n10380), .ZN(n10267) );
  NAND2_X1 U7862 ( .A1(n10520), .A2(n10267), .ZN(n10348) );
  INV_X1 U7863 ( .A(n10348), .ZN(n6607) );
  NOR2_X1 U7864 ( .A1(n10342), .A2(n6607), .ZN(n10241) );
  NAND2_X1 U7865 ( .A1(n8120), .A2(n6890), .ZN(n6609) );
  INV_X1 U7866 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8125) );
  OR2_X1 U7867 ( .A1(n5092), .A2(n8125), .ZN(n6608) );
  NAND2_X1 U7868 ( .A1(n6951), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6614) );
  OR2_X1 U7869 ( .A1(n6618), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6610) );
  AND2_X1 U7870 ( .A1(n6610), .A2(n6628), .ZN(n10394) );
  NAND2_X1 U7871 ( .A1(n6956), .A2(n10394), .ZN(n6613) );
  NAND2_X1 U7872 ( .A1(n6794), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6612) );
  NAND2_X1 U7873 ( .A1(n6898), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6611) );
  NAND2_X1 U7874 ( .A1(n8106), .A2(n6890), .ZN(n6616) );
  OR2_X1 U7875 ( .A1(n6692), .A2(n8084), .ZN(n6615) );
  NAND2_X1 U7876 ( .A1(n6951), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6622) );
  NAND2_X1 U7877 ( .A1(n6794), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6621) );
  NOR2_X1 U7878 ( .A1(n6637), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6617) );
  NOR2_X1 U7879 ( .A1(n6618), .A2(n6617), .ZN(n10405) );
  NAND2_X1 U7880 ( .A1(n6956), .A2(n10405), .ZN(n6620) );
  NAND2_X1 U7881 ( .A1(n6898), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6619) );
  NAND2_X1 U7882 ( .A1(n10537), .A2(n10262), .ZN(n10236) );
  INV_X1 U7883 ( .A(n10236), .ZN(n6623) );
  NAND2_X1 U7884 ( .A1(n7044), .A2(n6623), .ZN(n6624) );
  NAND2_X1 U7885 ( .A1(n10531), .A2(n10263), .ZN(n10237) );
  AND2_X1 U7886 ( .A1(n6624), .A2(n10237), .ZN(n6633) );
  NAND2_X1 U7887 ( .A1(n8261), .A2(n6890), .ZN(n6626) );
  OR2_X1 U7888 ( .A1(n6692), .A2(n9156), .ZN(n6625) );
  NAND2_X1 U7889 ( .A1(n6898), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U7890 ( .A1(n6951), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6631) );
  AOI21_X1 U7891 ( .B1(n10051), .B2(n6628), .A(n6627), .ZN(n10374) );
  NAND2_X1 U7892 ( .A1(n6956), .A2(n10374), .ZN(n6630) );
  NAND2_X1 U7893 ( .A1(n6794), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6629) );
  NAND2_X1 U7894 ( .A1(n10525), .A2(n10264), .ZN(n10238) );
  AND2_X1 U7895 ( .A1(n6633), .A2(n10238), .ZN(n7026) );
  INV_X1 U7896 ( .A(n7026), .ZN(n6919) );
  OR2_X1 U7897 ( .A1(n10537), .A2(n10262), .ZN(n7045) );
  NAND2_X1 U7898 ( .A1(n8040), .A2(n6890), .ZN(n6635) );
  AOI22_X1 U7899 ( .A1(n6895), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7950), .B2(
        n6894), .ZN(n6634) );
  NAND2_X1 U7900 ( .A1(n6898), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U7901 ( .A1(n6951), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6640) );
  NOR2_X1 U7902 ( .A1(n6902), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6636) );
  OR2_X1 U7903 ( .A1(n6637), .A2(n6636), .ZN(n10423) );
  INV_X1 U7904 ( .A(n10423), .ZN(n9943) );
  NAND2_X1 U7905 ( .A1(n6956), .A2(n9943), .ZN(n6639) );
  NAND2_X1 U7906 ( .A1(n6794), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6638) );
  OR2_X1 U7907 ( .A1(n10428), .A2(n10433), .ZN(n7025) );
  NAND2_X1 U7908 ( .A1(n7045), .A2(n7025), .ZN(n6643) );
  NAND2_X1 U7909 ( .A1(n10428), .A2(n10433), .ZN(n7111) );
  NAND2_X1 U7910 ( .A1(n10236), .A2(n7111), .ZN(n6642) );
  MUX2_X1 U7911 ( .A(n6643), .B(n6642), .S(n7547), .Z(n6644) );
  INV_X1 U7912 ( .A(n6644), .ZN(n6916) );
  NAND2_X1 U7913 ( .A1(n5731), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U7914 ( .A1(n6668), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6646) );
  NAND2_X1 U7915 ( .A1(n6681), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6645) );
  INV_X1 U7916 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7377) );
  OR2_X1 U7917 ( .A1(n7410), .A2(n7562), .ZN(n6649) );
  NAND2_X1 U7918 ( .A1(n6667), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6653) );
  NAND2_X1 U7919 ( .A1(n6681), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6652) );
  NAND2_X1 U7920 ( .A1(n5731), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6651) );
  NAND2_X1 U7921 ( .A1(n6668), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6650) );
  INV_X1 U7922 ( .A(SI_0_), .ZN(n6655) );
  INV_X1 U7923 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6654) );
  OAI21_X1 U7924 ( .B1(n7362), .B2(n6655), .A(n6654), .ZN(n6656) );
  AND2_X1 U7925 ( .A1(n6657), .A2(n6656), .ZN(n10587) );
  NAND2_X1 U7926 ( .A1(n7969), .A2(n7970), .ZN(n6659) );
  INV_X1 U7927 ( .A(n7077), .ZN(n8799) );
  INV_X1 U7928 ( .A(n10776), .ZN(n7981) );
  NAND2_X1 U7929 ( .A1(n8799), .A2(n7981), .ZN(n6658) );
  NAND2_X1 U7930 ( .A1(n6659), .A2(n6658), .ZN(n6745) );
  NAND2_X1 U7931 ( .A1(n6667), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U7932 ( .A1(n5091), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6662) );
  NAND2_X1 U7933 ( .A1(n5731), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6661) );
  NAND2_X1 U7934 ( .A1(n6681), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6660) );
  AND4_X2 U7935 ( .A1(n6663), .A2(n6662), .A3(n6661), .A4(n6660), .ZN(n7657)
         );
  OR2_X1 U7936 ( .A1(n6664), .A2(n6838), .ZN(n6673) );
  XNOR2_X1 U7937 ( .A(n6673), .B(P1_IR_REG_2__SCAN_IN), .ZN(n10745) );
  INV_X1 U7938 ( .A(n10745), .ZN(n7563) );
  INV_X1 U7939 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7360) );
  OR2_X1 U7940 ( .A1(n6676), .A2(n7364), .ZN(n6665) );
  OAI211_X1 U7941 ( .C1(n7410), .C2(n7563), .A(n6666), .B(n6665), .ZN(n7797)
         );
  INV_X1 U7942 ( .A(n7797), .ZN(n7799) );
  NAND2_X1 U7943 ( .A1(n6667), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6672) );
  NAND2_X1 U7944 ( .A1(n6668), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6670) );
  INV_X1 U7945 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8033) );
  NAND2_X1 U7946 ( .A1(n6681), .A2(n8033), .ZN(n6669) );
  INV_X1 U7947 ( .A(n8798), .ZN(n10103) );
  INV_X1 U7948 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9189) );
  NAND2_X1 U7949 ( .A1(n6673), .A2(n9189), .ZN(n6674) );
  NAND2_X1 U7950 ( .A1(n6674), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6675) );
  XNOR2_X1 U7951 ( .A(n6675), .B(P1_IR_REG_3__SCAN_IN), .ZN(n7595) );
  INV_X1 U7952 ( .A(n7595), .ZN(n7383) );
  INV_X1 U7953 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7385) );
  OR2_X1 U7954 ( .A1(n6676), .A2(n7384), .ZN(n6677) );
  OAI211_X1 U7955 ( .C1(n7410), .C2(n7383), .A(n6678), .B(n6677), .ZN(n8034)
         );
  NAND2_X1 U7956 ( .A1(n10103), .A2(n7806), .ZN(n7000) );
  AND2_X1 U7957 ( .A1(n7000), .A2(n6679), .ZN(n7082) );
  OAI21_X1 U7958 ( .B1(n6745), .B2(n10783), .A(n7082), .ZN(n6696) );
  NAND2_X1 U7959 ( .A1(n8798), .A2(n8034), .ZN(n7084) );
  NAND2_X1 U7960 ( .A1(n6667), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6686) );
  NAND2_X1 U7961 ( .A1(n6853), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6685) );
  NOR2_X1 U7962 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6680) );
  NOR2_X1 U7963 ( .A1(n6720), .A2(n6680), .ZN(n10828) );
  NAND2_X1 U7964 ( .A1(n6681), .A2(n10828), .ZN(n6684) );
  NAND2_X1 U7965 ( .A1(n5091), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6683) );
  INV_X1 U7966 ( .A(n8015), .ZN(n10102) );
  NAND2_X1 U7967 ( .A1(n6687), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6688) );
  MUX2_X1 U7968 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6688), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n6691) );
  NAND2_X1 U7969 ( .A1(n6691), .A2(n6690), .ZN(n7572) );
  OR2_X1 U7970 ( .A1(n6676), .A2(n7378), .ZN(n6694) );
  INV_X1 U7971 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7379) );
  OR2_X1 U7972 ( .A1(n6692), .A2(n7379), .ZN(n6693) );
  OAI211_X1 U7973 ( .C1(n7410), .C2(n7572), .A(n6694), .B(n6693), .ZN(n10829)
         );
  INV_X1 U7974 ( .A(n7046), .ZN(n6695) );
  AOI21_X1 U7975 ( .B1(n6696), .B2(n7084), .A(n6695), .ZN(n6730) );
  NAND2_X1 U7976 ( .A1(n6898), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6703) );
  NAND2_X1 U7977 ( .A1(n6853), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6702) );
  INV_X1 U7978 ( .A(n6719), .ZN(n6697) );
  AOI21_X1 U7979 ( .B1(n6697), .B2(P1_REG3_REG_6__SCAN_IN), .A(
        P1_REG3_REG_7__SCAN_IN), .ZN(n6698) );
  OR2_X1 U7980 ( .A1(n6698), .A2(n6731), .ZN(n8190) );
  INV_X1 U7981 ( .A(n8190), .ZN(n6699) );
  NAND2_X1 U7982 ( .A1(n6956), .A2(n6699), .ZN(n6701) );
  NAND2_X1 U7983 ( .A1(n6794), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6700) );
  NAND4_X1 U7984 ( .A1(n6703), .A2(n6702), .A3(n6701), .A4(n6700), .ZN(n10099)
         );
  INV_X1 U7985 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9187) );
  OR2_X1 U7986 ( .A1(n6692), .A2(n9187), .ZN(n6707) );
  NOR2_X1 U7987 ( .A1(n6690), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n6738) );
  OR2_X1 U7988 ( .A1(n6738), .A2(n6838), .ZN(n6713) );
  INV_X1 U7989 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8984) );
  NAND2_X1 U7990 ( .A1(n6713), .A2(n8984), .ZN(n6715) );
  NAND2_X1 U7991 ( .A1(n6715), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6705) );
  INV_X1 U7992 ( .A(n7706), .ZN(n7387) );
  OR2_X1 U7993 ( .A1(n7410), .A2(n7387), .ZN(n6706) );
  NAND2_X1 U7994 ( .A1(n6898), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6712) );
  NAND2_X1 U7995 ( .A1(n6853), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6711) );
  XNOR2_X1 U7996 ( .A(n6719), .B(P1_REG3_REG_6__SCAN_IN), .ZN(n8166) );
  NAND2_X1 U7997 ( .A1(n6956), .A2(n8166), .ZN(n6710) );
  NAND2_X1 U7998 ( .A1(n6794), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6709) );
  INV_X1 U7999 ( .A(n6713), .ZN(n6714) );
  NAND2_X1 U8000 ( .A1(n6714), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6716) );
  INV_X1 U8001 ( .A(n7620), .ZN(n7567) );
  OR2_X1 U8002 ( .A1(n6676), .A2(n7375), .ZN(n6718) );
  INV_X1 U8003 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7373) );
  OR2_X1 U8004 ( .A1(n6692), .A2(n7373), .ZN(n6717) );
  OAI211_X1 U8005 ( .C1(n7410), .C2(n7567), .A(n6718), .B(n6717), .ZN(n8149)
         );
  NAND2_X1 U8006 ( .A1(n8181), .A2(n8149), .ZN(n7987) );
  NAND2_X1 U8007 ( .A1(n8015), .A2(n10829), .ZN(n8011) );
  NAND2_X1 U8008 ( .A1(n6853), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U8009 ( .A1(n6794), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6724) );
  OAI21_X1 U8010 ( .B1(n6720), .B2(P1_REG3_REG_5__SCAN_IN), .A(n6719), .ZN(
        n6721) );
  INV_X1 U8011 ( .A(n6721), .ZN(n8079) );
  NAND2_X1 U8012 ( .A1(n6956), .A2(n8079), .ZN(n6723) );
  NAND2_X1 U8013 ( .A1(n6898), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6722) );
  AND4_X2 U8014 ( .A1(n6725), .A2(n6724), .A3(n6723), .A4(n6722), .ZN(n8071)
         );
  NAND2_X1 U8015 ( .A1(n6690), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6726) );
  XNOR2_X1 U8016 ( .A(n6726), .B(P1_IR_REG_5__SCAN_IN), .ZN(n7608) );
  INV_X1 U8017 ( .A(n7608), .ZN(n7380) );
  OR2_X1 U8018 ( .A1(n6676), .A2(n7381), .ZN(n6728) );
  INV_X1 U8019 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7382) );
  OR2_X1 U8020 ( .A1(n6692), .A2(n7382), .ZN(n6727) );
  OAI211_X1 U8021 ( .C1(n7410), .C2(n7380), .A(n6728), .B(n6727), .ZN(n8072)
         );
  NAND2_X1 U8022 ( .A1(n8071), .A2(n8072), .ZN(n7049) );
  NAND4_X1 U8023 ( .A1(n7987), .A2(n8011), .A3(n7049), .A4(n6976), .ZN(n6729)
         );
  OR3_X1 U8024 ( .A1(n6730), .A2(n8272), .A3(n6729), .ZN(n6756) );
  NAND2_X1 U8025 ( .A1(n6853), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6736) );
  NAND2_X1 U8026 ( .A1(n6898), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6735) );
  OR2_X1 U8027 ( .A1(n6731), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6732) );
  AND2_X1 U8028 ( .A1(n6773), .A2(n6732), .ZN(n10898) );
  NAND2_X1 U8029 ( .A1(n6956), .A2(n10898), .ZN(n6734) );
  NAND2_X1 U8030 ( .A1(n6794), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6733) );
  NAND2_X1 U8031 ( .A1(n6890), .A2(n7391), .ZN(n6743) );
  NOR2_X1 U8032 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n6737) );
  NAND2_X1 U8033 ( .A1(n6738), .A2(n6737), .ZN(n6740) );
  NAND2_X1 U8034 ( .A1(n6740), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6739) );
  MUX2_X1 U8035 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6739), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n6741) );
  INV_X1 U8036 ( .A(n7873), .ZN(n7394) );
  OR2_X1 U8037 ( .A1(n7410), .A2(n7394), .ZN(n6742) );
  OAI211_X1 U8038 ( .C1(n6692), .C2(n7396), .A(n6743), .B(n6742), .ZN(n10899)
         );
  NAND2_X1 U8039 ( .A1(n8303), .A2(n10899), .ZN(n8275) );
  INV_X1 U8040 ( .A(n10858), .ZN(n8192) );
  NAND2_X1 U8041 ( .A1(n5344), .A2(n8192), .ZN(n10882) );
  NAND2_X1 U8042 ( .A1(n8275), .A2(n10882), .ZN(n10885) );
  NAND2_X1 U8043 ( .A1(n8275), .A2(n6976), .ZN(n6783) );
  INV_X1 U8044 ( .A(n8303), .ZN(n10098) );
  INV_X1 U8045 ( .A(n10899), .ZN(n10881) );
  NAND2_X1 U8046 ( .A1(n10098), .A2(n10881), .ZN(n10884) );
  NAND2_X1 U8047 ( .A1(n10099), .A2(n10858), .ZN(n6744) );
  NAND2_X1 U8048 ( .A1(n10884), .A2(n6744), .ZN(n7005) );
  NAND2_X1 U8049 ( .A1(n10884), .A2(n7547), .ZN(n6757) );
  AOI22_X1 U8050 ( .A1(n10885), .A2(n6783), .B1(n7005), .B2(n6757), .ZN(n6755)
         );
  INV_X1 U8051 ( .A(n10783), .ZN(n10788) );
  NAND2_X1 U8052 ( .A1(n6745), .A2(n10788), .ZN(n6999) );
  NAND3_X1 U8053 ( .A1(n6999), .A2(n7084), .A3(n7081), .ZN(n6748) );
  INV_X1 U8054 ( .A(n8071), .ZN(n10101) );
  NAND4_X1 U8055 ( .A1(n7000), .A2(n7046), .A3(n7086), .A4(n7547), .ZN(n6746)
         );
  INV_X1 U8056 ( .A(n8181), .ZN(n10100) );
  NAND2_X1 U8057 ( .A1(n10100), .A2(n8002), .ZN(n7986) );
  NOR2_X1 U8058 ( .A1(n6746), .A2(n5536), .ZN(n6747) );
  NAND2_X1 U8059 ( .A1(n8011), .A2(n7049), .ZN(n6749) );
  NAND2_X1 U8060 ( .A1(n6749), .A2(n7086), .ZN(n7088) );
  NAND3_X1 U8061 ( .A1(n7088), .A2(n7547), .A3(n7987), .ZN(n6754) );
  NAND3_X1 U8062 ( .A1(n7986), .A2(n7086), .A3(n6976), .ZN(n6750) );
  OAI21_X1 U8063 ( .B1(n6976), .B2(n7986), .A(n6750), .ZN(n6751) );
  INV_X1 U8064 ( .A(n6751), .ZN(n6753) );
  OR2_X1 U8065 ( .A1(n7987), .A2(n7547), .ZN(n6752) );
  INV_X1 U8066 ( .A(n6757), .ZN(n6769) );
  NAND2_X1 U8067 ( .A1(n7400), .A2(n6890), .ZN(n6762) );
  NAND2_X1 U8068 ( .A1(n6808), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6780) );
  INV_X1 U8069 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6806) );
  NAND2_X1 U8070 ( .A1(n6780), .A2(n6806), .ZN(n6758) );
  NAND2_X1 U8071 ( .A1(n6758), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6759) );
  INV_X1 U8072 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6805) );
  NAND2_X1 U8073 ( .A1(n6759), .A2(n6805), .ZN(n6787) );
  OR2_X1 U8074 ( .A1(n6759), .A2(n6805), .ZN(n6760) );
  AOI22_X1 U8075 ( .A1(n6895), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6894), .B2(
        n10105), .ZN(n6761) );
  NAND2_X1 U8076 ( .A1(n6898), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6768) );
  NAND2_X1 U8077 ( .A1(n6853), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6767) );
  AND2_X1 U8078 ( .A1(n6775), .A2(n6763), .ZN(n6764) );
  NOR2_X1 U8079 ( .A1(n6791), .A2(n6764), .ZN(n8375) );
  NAND2_X1 U8080 ( .A1(n6956), .A2(n8375), .ZN(n6766) );
  NAND2_X1 U8081 ( .A1(n6794), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6765) );
  NAND4_X1 U8082 ( .A1(n6768), .A2(n6767), .A3(n6766), .A4(n6765), .ZN(n10096)
         );
  NAND2_X1 U8083 ( .A1(n10917), .A2(n10096), .ZN(n7096) );
  NAND2_X1 U8084 ( .A1(n6769), .A2(n7096), .ZN(n6771) );
  INV_X1 U8085 ( .A(n10096), .ZN(n8427) );
  INV_X1 U8086 ( .A(n10917), .ZN(n8583) );
  NAND2_X1 U8087 ( .A1(n7008), .A2(n6976), .ZN(n6770) );
  NAND2_X1 U8088 ( .A1(n6771), .A2(n6770), .ZN(n6785) );
  NAND2_X1 U8089 ( .A1(n6853), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6779) );
  NAND2_X1 U8090 ( .A1(n6898), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U8091 ( .A1(n6773), .A2(n6772), .ZN(n6774) );
  AND2_X1 U8092 ( .A1(n6775), .A2(n6774), .ZN(n8337) );
  NAND2_X1 U8093 ( .A1(n6956), .A2(n8337), .ZN(n6777) );
  NAND2_X1 U8094 ( .A1(n6794), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6776) );
  NAND2_X1 U8095 ( .A1(n7398), .A2(n6890), .ZN(n6782) );
  XNOR2_X1 U8096 ( .A(n6780), .B(P1_IR_REG_9__SCAN_IN), .ZN(n8220) );
  AOI22_X1 U8097 ( .A1(n6895), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6894), .B2(
        n8220), .ZN(n6781) );
  NAND2_X1 U8098 ( .A1(n6782), .A2(n6781), .ZN(n8345) );
  NAND2_X1 U8099 ( .A1(n8372), .A2(n8345), .ZN(n8277) );
  INV_X1 U8100 ( .A(n8277), .ZN(n6801) );
  INV_X1 U8101 ( .A(n8372), .ZN(n10097) );
  INV_X1 U8102 ( .A(n8345), .ZN(n10908) );
  NAND2_X1 U8103 ( .A1(n10097), .A2(n10908), .ZN(n8276) );
  INV_X1 U8104 ( .A(n8276), .ZN(n7004) );
  OAI22_X1 U8105 ( .A1(n6801), .A2(n6783), .B1(n6976), .B2(n7004), .ZN(n6784)
         );
  NAND3_X1 U8106 ( .A1(n6786), .A2(n6785), .A3(n6784), .ZN(n6821) );
  INV_X1 U8107 ( .A(n7008), .ZN(n6799) );
  NAND2_X1 U8108 ( .A1(n7416), .A2(n6890), .ZN(n6790) );
  NAND2_X1 U8109 ( .A1(n6787), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6788) );
  XNOR2_X1 U8110 ( .A(n6788), .B(P1_IR_REG_11__SCAN_IN), .ZN(n8390) );
  AOI22_X1 U8111 ( .A1(n6895), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6894), .B2(
        n8390), .ZN(n6789) );
  NAND2_X1 U8112 ( .A1(n6898), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6798) );
  NAND2_X1 U8113 ( .A1(n6853), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6797) );
  NOR2_X1 U8114 ( .A1(n6791), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6792) );
  OR2_X1 U8115 ( .A1(n6812), .A2(n6792), .ZN(n8617) );
  INV_X1 U8116 ( .A(n8617), .ZN(n6793) );
  NAND2_X1 U8117 ( .A1(n6956), .A2(n6793), .ZN(n6796) );
  NAND2_X1 U8118 ( .A1(n6794), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6795) );
  OAI211_X1 U8119 ( .C1(n6799), .C2(n8276), .A(n10939), .B(n7096), .ZN(n6800)
         );
  INV_X1 U8120 ( .A(n6800), .ZN(n6804) );
  NAND2_X1 U8121 ( .A1(n8619), .A2(n8746), .ZN(n7010) );
  NAND2_X1 U8122 ( .A1(n7010), .A2(n7008), .ZN(n7095) );
  AND2_X1 U8123 ( .A1(n6801), .A2(n7096), .ZN(n6802) );
  NOR2_X1 U8124 ( .A1(n7095), .A2(n6802), .ZN(n6803) );
  MUX2_X1 U8125 ( .A(n6804), .B(n6803), .S(n7547), .Z(n6820) );
  NAND2_X1 U8126 ( .A1(n7430), .A2(n6890), .ZN(n6811) );
  INV_X1 U8127 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8994) );
  NAND3_X1 U8128 ( .A1(n6806), .A2(n8994), .A3(n6805), .ZN(n6807) );
  OAI21_X1 U8129 ( .B1(n6808), .B2(n6807), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6809) );
  XNOR2_X1 U8130 ( .A(n6809), .B(P1_IR_REG_12__SCAN_IN), .ZN(n8594) );
  AOI22_X1 U8131 ( .A1(n6895), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6894), .B2(
        n8594), .ZN(n6810) );
  NAND2_X1 U8132 ( .A1(n6853), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6817) );
  NAND2_X1 U8133 ( .A1(n6794), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6816) );
  OR2_X1 U8134 ( .A1(n6812), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6813) );
  AND2_X1 U8135 ( .A1(n6829), .A2(n6813), .ZN(n10954) );
  NAND2_X1 U8136 ( .A1(n6956), .A2(n10954), .ZN(n6815) );
  NAND2_X1 U8137 ( .A1(n6898), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6814) );
  NAND2_X1 U8138 ( .A1(n10957), .A2(n10094), .ZN(n7011) );
  NAND2_X1 U8139 ( .A1(n7011), .A2(n7010), .ZN(n6818) );
  NAND2_X1 U8140 ( .A1(n8548), .A2(n10939), .ZN(n7099) );
  MUX2_X1 U8141 ( .A(n6818), .B(n7099), .S(n7547), .Z(n6819) );
  INV_X1 U8142 ( .A(n6863), .ZN(n6835) );
  NAND2_X1 U8143 ( .A1(n7471), .A2(n6890), .ZN(n6827) );
  NOR2_X1 U8144 ( .A1(n6822), .A2(n6838), .ZN(n6823) );
  MUX2_X1 U8145 ( .A(n6838), .B(n6823), .S(P1_IR_REG_13__SCAN_IN), .Z(n6825)
         );
  OR2_X1 U8146 ( .A1(n6825), .A2(n6824), .ZN(n10129) );
  AOI22_X1 U8147 ( .A1(n6895), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6894), .B2(
        n10124), .ZN(n6826) );
  NAND2_X1 U8148 ( .A1(n6853), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6834) );
  NAND2_X1 U8149 ( .A1(n6898), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6833) );
  NAND2_X1 U8150 ( .A1(n6829), .A2(n6828), .ZN(n6830) );
  AND2_X1 U8151 ( .A1(n6844), .A2(n6830), .ZN(n10044) );
  NAND2_X1 U8152 ( .A1(n6956), .A2(n10044), .ZN(n6832) );
  NAND2_X1 U8153 ( .A1(n6794), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6831) );
  OR2_X1 U8154 ( .A1(n9799), .A2(n9924), .ZN(n7012) );
  NAND3_X1 U8155 ( .A1(n6835), .A2(n7012), .A3(n8548), .ZN(n6836) );
  NAND2_X1 U8156 ( .A1(n9799), .A2(n9924), .ZN(n7015) );
  NAND2_X1 U8157 ( .A1(n6836), .A2(n7015), .ZN(n6861) );
  NAND2_X1 U8158 ( .A1(n7556), .A2(n6890), .ZN(n6842) );
  NOR2_X1 U8159 ( .A1(n6824), .A2(n6838), .ZN(n6837) );
  MUX2_X1 U8160 ( .A(n6838), .B(n6837), .S(P1_IR_REG_14__SCAN_IN), .Z(n6840)
         );
  INV_X1 U8161 ( .A(n6542), .ZN(n6839) );
  INV_X1 U8162 ( .A(n10131), .ZN(n10143) );
  AOI22_X1 U8163 ( .A1(n6895), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6894), .B2(
        n10143), .ZN(n6841) );
  NAND2_X1 U8164 ( .A1(n6898), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6849) );
  NAND2_X1 U8165 ( .A1(n6853), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6848) );
  NAND2_X1 U8166 ( .A1(n6844), .A2(n6843), .ZN(n6845) );
  AND2_X1 U8167 ( .A1(n6855), .A2(n6845), .ZN(n9922) );
  NAND2_X1 U8168 ( .A1(n6956), .A2(n9922), .ZN(n6847) );
  NAND2_X1 U8169 ( .A1(n6794), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6846) );
  NAND4_X1 U8170 ( .A1(n6849), .A2(n6848), .A3(n6847), .A4(n6846), .ZN(n10551)
         );
  INV_X1 U8171 ( .A(n10551), .ZN(n10257) );
  OR2_X1 U8172 ( .A1(n10255), .A2(n10257), .ZN(n7058) );
  NAND2_X1 U8173 ( .A1(n7642), .A2(n6890), .ZN(n6852) );
  XNOR2_X1 U8174 ( .A(n6850), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10158) );
  AOI22_X1 U8175 ( .A1(n6895), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6894), .B2(
        n10158), .ZN(n6851) );
  NAND2_X1 U8176 ( .A1(n6853), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6860) );
  NAND2_X1 U8177 ( .A1(n6794), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6859) );
  AND2_X1 U8178 ( .A1(n6855), .A2(n6854), .ZN(n6856) );
  NOR2_X1 U8179 ( .A1(n6870), .A2(n6856), .ZN(n10993) );
  NAND2_X1 U8180 ( .A1(n6956), .A2(n10993), .ZN(n6858) );
  NAND2_X1 U8181 ( .A1(n6898), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6857) );
  NAND2_X1 U8182 ( .A1(n10556), .A2(n10465), .ZN(n7016) );
  NAND2_X1 U8183 ( .A1(n10255), .A2(n10257), .ZN(n7057) );
  NAND2_X1 U8184 ( .A1(n7016), .A2(n7057), .ZN(n7101) );
  AND2_X1 U8185 ( .A1(n7015), .A2(n7011), .ZN(n7098) );
  INV_X1 U8186 ( .A(n7098), .ZN(n6862) );
  AND2_X1 U8187 ( .A1(n7058), .A2(n7012), .ZN(n7102) );
  OAI21_X1 U8188 ( .B1(n6863), .B2(n6862), .A(n7102), .ZN(n6865) );
  INV_X1 U8189 ( .A(n7018), .ZN(n6864) );
  NAND2_X1 U8190 ( .A1(n7689), .A2(n6890), .ZN(n6869) );
  XNOR2_X1 U8191 ( .A(n6867), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10182) );
  AOI22_X1 U8192 ( .A1(n6895), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6894), .B2(
        n10182), .ZN(n6868) );
  NAND2_X1 U8193 ( .A1(n6898), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6875) );
  NAND2_X1 U8194 ( .A1(n6853), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6874) );
  OR2_X1 U8195 ( .A1(n6870), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6871) );
  AND2_X1 U8196 ( .A1(n6871), .A2(n6882), .ZN(n10001) );
  NAND2_X1 U8197 ( .A1(n6956), .A2(n10001), .ZN(n6873) );
  NAND2_X1 U8198 ( .A1(n6794), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6872) );
  NAND2_X1 U8199 ( .A1(n10480), .A2(n10450), .ZN(n7104) );
  NAND2_X1 U8200 ( .A1(n7104), .A2(n7016), .ZN(n6876) );
  OR2_X1 U8201 ( .A1(n10480), .A2(n10450), .ZN(n7020) );
  NAND2_X1 U8202 ( .A1(n7020), .A2(n7018), .ZN(n7106) );
  MUX2_X1 U8203 ( .A(n6876), .B(n7106), .S(n6976), .Z(n6889) );
  NAND2_X1 U8204 ( .A1(n7817), .A2(n6890), .ZN(n6880) );
  NAND2_X1 U8205 ( .A1(n6867), .A2(n9211), .ZN(n6877) );
  NAND2_X1 U8206 ( .A1(n6877), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6878) );
  XNOR2_X1 U8207 ( .A(n6878), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10198) );
  AOI22_X1 U8208 ( .A1(n6895), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6894), .B2(
        n10198), .ZN(n6879) );
  NAND2_X1 U8209 ( .A1(n6898), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6887) );
  NAND2_X1 U8210 ( .A1(n6951), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6886) );
  NAND2_X1 U8211 ( .A1(n6882), .A2(n6881), .ZN(n6883) );
  AND2_X1 U8212 ( .A1(n6900), .A2(n6883), .ZN(n10453) );
  NAND2_X1 U8213 ( .A1(n6956), .A2(n10453), .ZN(n6885) );
  NAND2_X1 U8214 ( .A1(n6794), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6884) );
  NAND2_X1 U8215 ( .A1(n10543), .A2(n10463), .ZN(n7022) );
  NAND2_X1 U8216 ( .A1(n7107), .A2(n7022), .ZN(n10445) );
  INV_X1 U8217 ( .A(n10445), .ZN(n10447) );
  MUX2_X1 U8218 ( .A(n7104), .B(n7020), .S(n7547), .Z(n6888) );
  NAND2_X1 U8219 ( .A1(n7821), .A2(n6890), .ZN(n6897) );
  NAND2_X1 U8220 ( .A1(n6891), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n6892) );
  AND2_X1 U8221 ( .A1(n6893), .A2(n6892), .ZN(n10209) );
  AOI22_X1 U8222 ( .A1(n6895), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6894), .B2(
        n10209), .ZN(n6896) );
  NAND2_X1 U8223 ( .A1(n6898), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6906) );
  NAND2_X1 U8224 ( .A1(n6951), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6905) );
  AND2_X1 U8225 ( .A1(n6900), .A2(n6899), .ZN(n6901) );
  NOR2_X1 U8226 ( .A1(n6902), .A2(n6901), .ZN(n10439) );
  NAND2_X1 U8227 ( .A1(n6956), .A2(n10439), .ZN(n6904) );
  NAND2_X1 U8228 ( .A1(n6794), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6903) );
  NAND4_X1 U8229 ( .A1(n6906), .A2(n6905), .A3(n6904), .A4(n6903), .ZN(n10417)
         );
  OR2_X1 U8230 ( .A1(n10260), .A2(n10451), .ZN(n7024) );
  AND2_X1 U8231 ( .A1(n10260), .A2(n10451), .ZN(n7023) );
  INV_X1 U8232 ( .A(n7023), .ZN(n6907) );
  NAND3_X1 U8233 ( .A1(n6908), .A2(n7111), .A3(n6907), .ZN(n6914) );
  AND2_X1 U8234 ( .A1(n7025), .A2(n7024), .ZN(n7114) );
  INV_X1 U8235 ( .A(n7022), .ZN(n6909) );
  OR2_X1 U8236 ( .A1(n7023), .A2(n6909), .ZN(n7110) );
  INV_X1 U8237 ( .A(n7110), .ZN(n6910) );
  NAND2_X1 U8238 ( .A1(n6911), .A2(n6910), .ZN(n6912) );
  NAND2_X1 U8239 ( .A1(n7114), .A2(n6912), .ZN(n6913) );
  INV_X1 U8240 ( .A(n7044), .ZN(n6917) );
  NOR2_X1 U8241 ( .A1(n6921), .A2(n6917), .ZN(n6918) );
  NOR2_X1 U8242 ( .A1(n6919), .A2(n6918), .ZN(n6922) );
  NAND2_X1 U8243 ( .A1(n7044), .A2(n7045), .ZN(n7116) );
  INV_X1 U8244 ( .A(n7116), .ZN(n6920) );
  OR2_X1 U8245 ( .A1(n10525), .A2(n10264), .ZN(n7043) );
  OR2_X1 U8246 ( .A1(n10520), .A2(n10267), .ZN(n7042) );
  NAND2_X1 U8247 ( .A1(n7042), .A2(n7043), .ZN(n6993) );
  NAND2_X1 U8248 ( .A1(n10241), .A2(n6923), .ZN(n6933) );
  NAND2_X1 U8249 ( .A1(n8632), .A2(n6890), .ZN(n6925) );
  INV_X1 U8250 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8651) );
  OR2_X1 U8251 ( .A1(n6692), .A2(n8651), .ZN(n6924) );
  NAND2_X1 U8252 ( .A1(n6951), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6932) );
  NAND2_X1 U8253 ( .A1(n6898), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6931) );
  INV_X1 U8254 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6926) );
  NAND2_X1 U8255 ( .A1(n6927), .A2(n6926), .ZN(n6928) );
  AND2_X1 U8256 ( .A1(n6942), .A2(n6928), .ZN(n10331) );
  NAND2_X1 U8257 ( .A1(n6956), .A2(n10331), .ZN(n6930) );
  NAND2_X1 U8258 ( .A1(n5091), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6929) );
  NAND4_X1 U8259 ( .A1(n6932), .A2(n6931), .A3(n6930), .A4(n6929), .ZN(n10351)
         );
  OR2_X1 U8260 ( .A1(n10510), .A2(n10318), .ZN(n6997) );
  NAND2_X1 U8261 ( .A1(n10510), .A2(n10318), .ZN(n10242) );
  NAND3_X1 U8262 ( .A1(n6933), .A2(n10334), .A3(n10239), .ZN(n6938) );
  NAND2_X1 U8263 ( .A1(n10348), .A2(n10238), .ZN(n6934) );
  INV_X1 U8264 ( .A(n10342), .ZN(n10349) );
  OAI211_X1 U8265 ( .C1(n6935), .C2(n6934), .A(n10349), .B(n7042), .ZN(n6936)
         );
  NAND2_X1 U8266 ( .A1(n6936), .A2(n7027), .ZN(n6937) );
  NAND2_X1 U8267 ( .A1(n8779), .A2(n6890), .ZN(n6940) );
  OR2_X1 U8268 ( .A1(n6692), .A2(n9148), .ZN(n6939) );
  NAND2_X1 U8269 ( .A1(n6951), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6947) );
  NAND2_X1 U8270 ( .A1(n6898), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6946) );
  INV_X1 U8271 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6941) );
  NAND2_X1 U8272 ( .A1(n6942), .A2(n6941), .ZN(n6943) );
  AND2_X1 U8273 ( .A1(n6953), .A2(n6943), .ZN(n10323) );
  NAND2_X1 U8274 ( .A1(n6956), .A2(n10323), .ZN(n6945) );
  NAND2_X1 U8275 ( .A1(n5091), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6944) );
  NAND2_X1 U8276 ( .A1(n10506), .A2(n10305), .ZN(n7040) );
  INV_X1 U8277 ( .A(n7040), .ZN(n10243) );
  AND2_X1 U8278 ( .A1(n7040), .A2(n10242), .ZN(n7030) );
  INV_X1 U8279 ( .A(n7030), .ZN(n6948) );
  AND2_X1 U8280 ( .A1(n6948), .A2(n6976), .ZN(n6963) );
  NAND2_X1 U8281 ( .A1(n8755), .A2(n6890), .ZN(n6950) );
  OR2_X1 U8282 ( .A1(n5092), .A2(n9149), .ZN(n6949) );
  NAND2_X1 U8283 ( .A1(n6951), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6960) );
  NAND2_X1 U8284 ( .A1(n6898), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6959) );
  INV_X1 U8285 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6952) );
  NAND2_X1 U8286 ( .A1(n6953), .A2(n6952), .ZN(n6954) );
  NAND2_X1 U8287 ( .A1(n6956), .A2(n10308), .ZN(n6958) );
  NAND2_X1 U8288 ( .A1(n6794), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6957) );
  NAND2_X1 U8289 ( .A1(n10501), .A2(n10319), .ZN(n10245) );
  NOR2_X1 U8290 ( .A1(n7041), .A2(n7547), .ZN(n6961) );
  NOR2_X1 U8291 ( .A1(n10302), .A2(n6961), .ZN(n6962) );
  OAI21_X1 U8292 ( .B1(n6964), .B2(n6963), .A(n6962), .ZN(n6967) );
  NAND2_X1 U8293 ( .A1(n10495), .A2(n10306), .ZN(n10247) );
  NAND2_X1 U8294 ( .A1(n6965), .A2(n10247), .ZN(n10291) );
  INV_X1 U8295 ( .A(n10291), .ZN(n10283) );
  MUX2_X1 U8296 ( .A(n10245), .B(n6992), .S(n7547), .Z(n6966) );
  NAND3_X1 U8297 ( .A1(n6967), .A2(n10283), .A3(n6966), .ZN(n6970) );
  NAND2_X1 U8298 ( .A1(n7125), .A2(n10247), .ZN(n6968) );
  NAND2_X1 U8299 ( .A1(n6968), .A2(n7547), .ZN(n6969) );
  NAND3_X1 U8300 ( .A1(n6971), .A2(n6970), .A3(n6969), .ZN(n6972) );
  NAND3_X1 U8301 ( .A1(n7036), .A2(n6973), .A3(n6972), .ZN(n6975) );
  INV_X1 U8302 ( .A(n10250), .ZN(n10092) );
  NAND2_X1 U8303 ( .A1(n10092), .A2(n10091), .ZN(n6974) );
  NAND2_X1 U8304 ( .A1(n10226), .A2(n6974), .ZN(n7033) );
  MUX2_X1 U8305 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7362), .Z(n6980) );
  INV_X1 U8306 ( .A(SI_31_), .ZN(n9045) );
  XNOR2_X1 U8307 ( .A(n6980), .B(n9045), .ZN(n6981) );
  INV_X1 U8308 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10578) );
  NOR2_X1 U8309 ( .A1(n6692), .A2(n10578), .ZN(n6982) );
  AND2_X1 U8310 ( .A1(n10484), .A2(n10091), .ZN(n7037) );
  INV_X1 U8311 ( .A(n7037), .ZN(n7131) );
  NAND2_X1 U8312 ( .A1(n6983), .A2(n7131), .ZN(n6986) );
  INV_X1 U8313 ( .A(n10484), .ZN(n6984) );
  NAND2_X1 U8314 ( .A1(n6984), .A2(n10230), .ZN(n7130) );
  AOI21_X1 U8315 ( .B1(n7130), .B2(n7036), .A(n7547), .ZN(n6985) );
  AOI21_X1 U8316 ( .B1(n6986), .B2(n7130), .A(n6985), .ZN(n7144) );
  INV_X1 U8317 ( .A(n6988), .ZN(n6989) );
  NAND2_X1 U8318 ( .A1(n6989), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6990) );
  INV_X1 U8319 ( .A(n7525), .ZN(n7546) );
  NAND2_X1 U8320 ( .A1(n7161), .A2(n7546), .ZN(n7541) );
  INV_X1 U8321 ( .A(n7541), .ZN(n6991) );
  OAI211_X1 U8322 ( .C1(n7131), .C2(n10219), .A(n6991), .B(n5452), .ZN(n7143)
         );
  NAND2_X1 U8323 ( .A1(n6992), .A2(n7041), .ZN(n7031) );
  NAND2_X1 U8324 ( .A1(n6993), .A2(n10348), .ZN(n6994) );
  NAND2_X1 U8325 ( .A1(n10239), .A2(n6994), .ZN(n6995) );
  NAND2_X1 U8326 ( .A1(n6995), .A2(n7027), .ZN(n6996) );
  NAND2_X1 U8327 ( .A1(n6997), .A2(n6996), .ZN(n6998) );
  NOR2_X1 U8328 ( .A1(n7031), .A2(n6998), .ZN(n7074) );
  NAND2_X1 U8329 ( .A1(n6999), .A2(n7081), .ZN(n8028) );
  INV_X1 U8330 ( .A(n8032), .ZN(n7001) );
  NAND2_X1 U8331 ( .A1(n8028), .A2(n7001), .ZN(n7002) );
  NAND2_X1 U8332 ( .A1(n7002), .A2(n7084), .ZN(n10817) );
  NAND2_X1 U8333 ( .A1(n10817), .A2(n7046), .ZN(n8012) );
  INV_X1 U8334 ( .A(n7086), .ZN(n7003) );
  NOR2_X1 U8335 ( .A1(n7005), .A2(n7004), .ZN(n7053) );
  NAND2_X1 U8336 ( .A1(n8184), .A2(n7053), .ZN(n7007) );
  NAND3_X1 U8337 ( .A1(n10885), .A2(n8276), .A3(n10884), .ZN(n7006) );
  AND2_X1 U8338 ( .A1(n7006), .A2(n8277), .ZN(n7093) );
  NAND2_X1 U8339 ( .A1(n7007), .A2(n7093), .ZN(n8365) );
  NAND2_X1 U8340 ( .A1(n7096), .A2(n7008), .ZN(n8425) );
  INV_X1 U8341 ( .A(n8425), .ZN(n8366) );
  NAND2_X1 U8342 ( .A1(n8365), .A2(n8366), .ZN(n7009) );
  NAND2_X1 U8343 ( .A1(n10939), .A2(n7010), .ZN(n8555) );
  NAND2_X1 U8344 ( .A1(n8548), .A2(n7011), .ZN(n10938) );
  INV_X1 U8345 ( .A(n10938), .ZN(n10940) );
  NAND2_X1 U8346 ( .A1(n7012), .A2(n7015), .ZN(n8635) );
  INV_X1 U8347 ( .A(n8548), .ZN(n7013) );
  NOR2_X1 U8348 ( .A1(n8635), .A2(n7013), .ZN(n7014) );
  NAND2_X1 U8349 ( .A1(n10946), .A2(n7014), .ZN(n8550) );
  INV_X1 U8350 ( .A(n10548), .ZN(n7017) );
  NAND2_X1 U8351 ( .A1(n7019), .A2(n7018), .ZN(n10459) );
  NAND2_X1 U8352 ( .A1(n7020), .A2(n7104), .ZN(n10469) );
  INV_X1 U8353 ( .A(n10469), .ZN(n7021) );
  AOI21_X2 U8354 ( .B1(n10432), .B2(n7024), .A(n7023), .ZN(n10416) );
  NAND2_X1 U8355 ( .A1(n7025), .A2(n7111), .ZN(n10419) );
  OAI21_X2 U8356 ( .B1(n10416), .B2(n10419), .A(n7111), .ZN(n10409) );
  INV_X1 U8357 ( .A(n10409), .ZN(n7029) );
  AND2_X1 U8358 ( .A1(n7026), .A2(n10348), .ZN(n7028) );
  AND2_X1 U8359 ( .A1(n7028), .A2(n7027), .ZN(n7075) );
  OAI21_X1 U8360 ( .B1(n7029), .B2(n7116), .A(n7075), .ZN(n7032) );
  OAI211_X1 U8361 ( .C1(n7031), .C2(n7030), .A(n10245), .B(n10247), .ZN(n7121)
         );
  AOI21_X1 U8362 ( .B1(n7074), .B2(n7032), .A(n7121), .ZN(n7034) );
  OAI211_X1 U8363 ( .C1(n7127), .C2(n7034), .A(n7125), .B(n7033), .ZN(n7035)
         );
  AOI21_X1 U8364 ( .B1(n7036), .B2(n7035), .A(n7037), .ZN(n7072) );
  NAND2_X1 U8365 ( .A1(n7130), .A2(n7656), .ZN(n7071) );
  AND2_X1 U8366 ( .A1(n10226), .A2(n10250), .ZN(n7123) );
  NOR2_X1 U8367 ( .A1(n7123), .A2(n7038), .ZN(n7070) );
  INV_X1 U8368 ( .A(n10315), .ZN(n10244) );
  NAND2_X1 U8369 ( .A1(n7043), .A2(n10238), .ZN(n10369) );
  INV_X1 U8370 ( .A(n10369), .ZN(n10379) );
  NAND2_X1 U8371 ( .A1(n7044), .A2(n10237), .ZN(n10391) );
  INV_X1 U8372 ( .A(n8635), .ZN(n7056) );
  NOR2_X1 U8373 ( .A1(n10818), .A2(n8032), .ZN(n7048) );
  AND2_X1 U8374 ( .A1(n7973), .A2(n7977), .ZN(n7076) );
  OR2_X1 U8375 ( .A1(n7076), .A2(n7970), .ZN(n7943) );
  NOR2_X1 U8376 ( .A1(n7943), .A2(n7161), .ZN(n7047) );
  AND4_X1 U8377 ( .A1(n7048), .A2(n7047), .A3(n10788), .A4(n7987), .ZN(n7052)
         );
  INV_X1 U8378 ( .A(n10885), .ZN(n7051) );
  NAND2_X1 U8379 ( .A1(n7049), .A2(n7086), .ZN(n8020) );
  NAND4_X1 U8380 ( .A1(n7052), .A2(n7051), .A3(n7050), .A4(n8277), .ZN(n7054)
         );
  NAND2_X1 U8381 ( .A1(n7053), .A2(n7986), .ZN(n7090) );
  NOR4_X1 U8382 ( .A1(n7054), .A2(n8555), .A3(n7090), .A4(n8425), .ZN(n7055)
         );
  NAND3_X1 U8383 ( .A1(n7056), .A2(n7055), .A3(n10940), .ZN(n7059) );
  NAND2_X1 U8384 ( .A1(n7058), .A2(n7057), .ZN(n8638) );
  NOR2_X1 U8385 ( .A1(n7059), .A2(n8638), .ZN(n7060) );
  NAND2_X1 U8386 ( .A1(n10548), .A2(n7060), .ZN(n7061) );
  NOR2_X1 U8387 ( .A1(n10469), .A2(n7061), .ZN(n7063) );
  XNOR2_X1 U8388 ( .A(n10260), .B(n10451), .ZN(n10436) );
  NOR2_X1 U8389 ( .A1(n10419), .A2(n10436), .ZN(n7062) );
  NAND4_X1 U8390 ( .A1(n10410), .A2(n10447), .A3(n7063), .A4(n7062), .ZN(n7064) );
  NOR2_X1 U8391 ( .A1(n10391), .A2(n7064), .ZN(n7065) );
  NAND3_X1 U8392 ( .A1(n10362), .A2(n10379), .A3(n7065), .ZN(n7066) );
  NOR2_X1 U8393 ( .A1(n10342), .A2(n7066), .ZN(n7067) );
  NAND3_X1 U8394 ( .A1(n10244), .A2(n10334), .A3(n7067), .ZN(n7068) );
  NOR2_X1 U8395 ( .A1(n10302), .A2(n7068), .ZN(n7069) );
  NAND4_X1 U8396 ( .A1(n7131), .A2(n7070), .A3(n7130), .A4(n5728), .ZN(n7135)
         );
  OAI21_X1 U8397 ( .B1(n7072), .B2(n7071), .A(n7135), .ZN(n7073) );
  INV_X1 U8398 ( .A(n7073), .ZN(n7137) );
  INV_X1 U8399 ( .A(n7074), .ZN(n7120) );
  INV_X1 U8400 ( .A(n7075), .ZN(n7118) );
  INV_X1 U8401 ( .A(n7076), .ZN(n7079) );
  NAND2_X1 U8402 ( .A1(n7077), .A2(n10776), .ZN(n7078) );
  NAND3_X1 U8403 ( .A1(n7079), .A2(n7161), .A3(n7078), .ZN(n7080) );
  NAND2_X1 U8404 ( .A1(n7081), .A2(n7080), .ZN(n7083) );
  OAI21_X1 U8405 ( .B1(n6745), .B2(n7083), .A(n7082), .ZN(n7085) );
  NAND2_X1 U8406 ( .A1(n7085), .A2(n7084), .ZN(n7087) );
  NAND3_X1 U8407 ( .A1(n7087), .A2(n7086), .A3(n7046), .ZN(n7089) );
  NAND3_X1 U8408 ( .A1(n7089), .A2(n7987), .A3(n7088), .ZN(n7092) );
  INV_X1 U8409 ( .A(n7090), .ZN(n7091) );
  NAND2_X1 U8410 ( .A1(n7092), .A2(n7091), .ZN(n7094) );
  NAND2_X1 U8411 ( .A1(n7094), .A2(n7093), .ZN(n7097) );
  AOI21_X1 U8412 ( .B1(n7097), .B2(n7096), .A(n7095), .ZN(n7100) );
  OAI21_X1 U8413 ( .B1(n7100), .B2(n7099), .A(n7098), .ZN(n7103) );
  AOI21_X1 U8414 ( .B1(n7103), .B2(n7102), .A(n7101), .ZN(n7105) );
  OAI21_X1 U8415 ( .B1(n7106), .B2(n7105), .A(n7104), .ZN(n7108) );
  AND2_X1 U8416 ( .A1(n7108), .A2(n7107), .ZN(n7109) );
  OR2_X1 U8417 ( .A1(n7110), .A2(n7109), .ZN(n7113) );
  INV_X1 U8418 ( .A(n7111), .ZN(n7112) );
  AOI21_X1 U8419 ( .B1(n7114), .B2(n7113), .A(n7112), .ZN(n7115) );
  NOR2_X1 U8420 ( .A1(n7116), .A2(n7115), .ZN(n7117) );
  NOR2_X1 U8421 ( .A1(n7118), .A2(n7117), .ZN(n7119) );
  NOR2_X1 U8422 ( .A1(n7120), .A2(n7119), .ZN(n7122) );
  NOR2_X1 U8423 ( .A1(n7122), .A2(n7121), .ZN(n7126) );
  INV_X1 U8424 ( .A(n7123), .ZN(n7124) );
  OAI211_X1 U8425 ( .C1(n7127), .C2(n7126), .A(n7125), .B(n7124), .ZN(n7128)
         );
  NAND3_X1 U8426 ( .A1(n7130), .A2(n7129), .A3(n7128), .ZN(n7132) );
  NAND2_X1 U8427 ( .A1(n7132), .A2(n7131), .ZN(n7149) );
  AOI21_X1 U8428 ( .B1(n7149), .B2(n7950), .A(n7546), .ZN(n7133) );
  INV_X1 U8429 ( .A(n7133), .ZN(n7136) );
  NAND2_X1 U8430 ( .A1(n7950), .A2(n7509), .ZN(n7542) );
  OAI21_X1 U8431 ( .B1(n7161), .B2(n10219), .A(n7542), .ZN(n7134) );
  NAND2_X1 U8432 ( .A1(n7135), .A2(n7134), .ZN(n7139) );
  INV_X1 U8433 ( .A(n7138), .ZN(n7142) );
  INV_X1 U8434 ( .A(n7139), .ZN(n7140) );
  OAI211_X1 U8435 ( .C1(n7144), .C2(n7143), .A(n7142), .B(n7141), .ZN(n7145)
         );
  NAND2_X1 U8436 ( .A1(n7146), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7147) );
  OR2_X1 U8437 ( .A1(n7809), .A2(P1_U3086), .ZN(n8419) );
  INV_X1 U8438 ( .A(n8419), .ZN(n7148) );
  INV_X1 U8439 ( .A(n7151), .ZN(n10228) );
  NAND2_X1 U8440 ( .A1(n10746), .A2(n10228), .ZN(n7568) );
  NAND2_X1 U8441 ( .A1(n7152), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7153) );
  MUX2_X1 U8442 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7153), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n7154) );
  NAND2_X1 U8443 ( .A1(n7158), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7159) );
  NOR2_X2 U8444 ( .A1(n8653), .A2(n8587), .ZN(n7160) );
  INV_X1 U8445 ( .A(n10573), .ZN(n7162) );
  NAND2_X1 U8446 ( .A1(n7507), .A2(n7509), .ZN(n7544) );
  NAND2_X1 U8447 ( .A1(n7161), .A2(n7525), .ZN(n7512) );
  OR2_X1 U8448 ( .A1(n7544), .A2(n7512), .ZN(n7543) );
  NOR3_X1 U8449 ( .A1(n7568), .A2(n7162), .A3(n7543), .ZN(n7164) );
  OAI21_X1 U8450 ( .B1(n8419), .B2(n7509), .A(P1_B_REG_SCAN_IN), .ZN(n7163) );
  OAI22_X1 U8451 ( .A1(n7166), .A2(n7165), .B1(n7164), .B2(n7163), .ZN(
        P1_U3242) );
  AOI21_X1 U8452 ( .B1(n5125), .B2(n7167), .A(n7306), .ZN(n7278) );
  OAI21_X1 U8453 ( .B1(n8820), .B2(n9611), .A(n7167), .ZN(n7170) );
  INV_X1 U8454 ( .A(n7168), .ZN(n7169) );
  MUX2_X1 U8455 ( .A(n7170), .B(n7169), .S(n7739), .Z(n7276) );
  NAND2_X1 U8456 ( .A1(n7267), .A2(n7258), .ZN(n7172) );
  NAND2_X1 U8457 ( .A1(n7268), .A2(n7265), .ZN(n7171) );
  MUX2_X1 U8458 ( .A(n7172), .B(n7171), .S(n7306), .Z(n7270) );
  AND2_X1 U8459 ( .A1(n7252), .A2(n7175), .ZN(n7173) );
  MUX2_X1 U8460 ( .A(n7249), .B(n7173), .S(n7306), .Z(n7251) );
  OAI211_X1 U8461 ( .C1(n8534), .C2(n7176), .A(n7175), .B(n7174), .ZN(n7177)
         );
  MUX2_X1 U8462 ( .A(n8622), .B(n7177), .S(n7739), .Z(n7178) );
  INV_X1 U8463 ( .A(n7178), .ZN(n7250) );
  AND2_X1 U8464 ( .A1(n7203), .A2(n7917), .ZN(n7214) );
  NAND2_X1 U8465 ( .A1(n7202), .A2(n7179), .ZN(n7181) );
  INV_X1 U8466 ( .A(n7201), .ZN(n7180) );
  AOI21_X1 U8467 ( .B1(n7214), .B2(n7181), .A(n7180), .ZN(n7208) );
  NAND2_X1 U8468 ( .A1(n9405), .A2(n7889), .ZN(n7182) );
  NAND2_X1 U8469 ( .A1(n7736), .A2(n7182), .ZN(n8356) );
  NAND2_X1 U8470 ( .A1(n7183), .A2(n7182), .ZN(n7184) );
  NAND2_X1 U8471 ( .A1(n7184), .A2(n7185), .ZN(n7187) );
  OAI21_X1 U8472 ( .B1(n8356), .B2(n7730), .A(n7187), .ZN(n7186) );
  NAND2_X1 U8473 ( .A1(n7186), .A2(n7185), .ZN(n7189) );
  INV_X1 U8474 ( .A(n7187), .ZN(n7188) );
  MUX2_X1 U8475 ( .A(n7189), .B(n7188), .S(n7739), .Z(n7190) );
  NAND2_X1 U8476 ( .A1(n7190), .A2(n7633), .ZN(n7197) );
  NAND2_X1 U8477 ( .A1(n7213), .A2(n7191), .ZN(n7194) );
  NAND2_X1 U8478 ( .A1(n7199), .A2(n7192), .ZN(n7193) );
  MUX2_X1 U8479 ( .A(n7194), .B(n7193), .S(n7739), .Z(n7195) );
  INV_X1 U8480 ( .A(n7195), .ZN(n7196) );
  NAND2_X1 U8481 ( .A1(n7197), .A2(n7196), .ZN(n7198) );
  NAND2_X1 U8482 ( .A1(n7198), .A2(n7682), .ZN(n7212) );
  OAI211_X1 U8483 ( .C1(n7212), .C2(n5486), .A(n7917), .B(n7200), .ZN(n7206)
         );
  AND2_X1 U8484 ( .A1(n7202), .A2(n7201), .ZN(n7205) );
  INV_X1 U8485 ( .A(n7203), .ZN(n7204) );
  AOI21_X1 U8486 ( .B1(n7206), .B2(n7205), .A(n7204), .ZN(n7207) );
  MUX2_X1 U8487 ( .A(n7208), .B(n7207), .S(n7306), .Z(n7217) );
  NAND3_X1 U8488 ( .A1(n7218), .A2(n7739), .A3(n7209), .ZN(n7211) );
  AND2_X1 U8489 ( .A1(n7224), .A2(n7306), .ZN(n7210) );
  NAND2_X1 U8490 ( .A1(n7225), .A2(n7210), .ZN(n7220) );
  NAND2_X1 U8491 ( .A1(n7211), .A2(n7220), .ZN(n7228) );
  INV_X1 U8492 ( .A(n7212), .ZN(n7215) );
  NAND4_X1 U8493 ( .A1(n7215), .A2(n7739), .A3(n7214), .A4(n7213), .ZN(n7216)
         );
  NAND4_X1 U8494 ( .A1(n7217), .A2(n6451), .A3(n7228), .A4(n7216), .ZN(n7233)
         );
  OAI21_X1 U8495 ( .B1(n7220), .B2(n7219), .A(n7218), .ZN(n7221) );
  NOR2_X1 U8496 ( .A1(n7222), .A2(n7221), .ZN(n7231) );
  NAND2_X1 U8497 ( .A1(n7224), .A2(n7223), .ZN(n7227) );
  INV_X1 U8498 ( .A(n7225), .ZN(n7226) );
  AOI21_X1 U8499 ( .B1(n7228), .B2(n7227), .A(n7226), .ZN(n7229) );
  AND2_X1 U8500 ( .A1(n7236), .A2(n7229), .ZN(n7230) );
  MUX2_X1 U8501 ( .A(n7231), .B(n7230), .S(n7739), .Z(n7232) );
  NAND2_X1 U8502 ( .A1(n7233), .A2(n7232), .ZN(n7245) );
  INV_X1 U8503 ( .A(n7234), .ZN(n7235) );
  NOR2_X1 U8504 ( .A1(n7236), .A2(n7235), .ZN(n7238) );
  NOR2_X1 U8505 ( .A1(n7239), .A2(n8266), .ZN(n7244) );
  MUX2_X1 U8506 ( .A(n7241), .B(n7240), .S(n7739), .Z(n7242) );
  NAND2_X1 U8507 ( .A1(n8461), .A2(n7242), .ZN(n7243) );
  AOI21_X1 U8508 ( .B1(n7245), .B2(n7244), .A(n7243), .ZN(n7247) );
  NOR2_X1 U8509 ( .A1(n8528), .A2(n7739), .ZN(n7246) );
  OAI21_X1 U8510 ( .B1(n7247), .B2(n7246), .A(n8529), .ZN(n7248) );
  MUX2_X1 U8511 ( .A(n7253), .B(n7252), .S(n7739), .Z(n7254) );
  MUX2_X1 U8512 ( .A(n9389), .B(n9321), .S(n7739), .Z(n7255) );
  NAND2_X1 U8513 ( .A1(n7256), .A2(n7255), .ZN(n7261) );
  NAND3_X1 U8514 ( .A1(n7261), .A2(n9321), .A3(n7264), .ZN(n7259) );
  NAND3_X1 U8515 ( .A1(n8699), .A2(n7262), .A3(n8809), .ZN(n7257) );
  NAND3_X1 U8516 ( .A1(n7261), .A2(n9389), .A3(n7260), .ZN(n7266) );
  INV_X1 U8517 ( .A(n9321), .ZN(n8727) );
  NAND3_X1 U8518 ( .A1(n8699), .A2(n7262), .A3(n8727), .ZN(n7263) );
  MUX2_X1 U8519 ( .A(n7268), .B(n7267), .S(n7306), .Z(n7269) );
  MUX2_X1 U8520 ( .A(n7272), .B(n7271), .S(n7306), .Z(n7273) );
  AND3_X1 U8521 ( .A1(n9627), .A2(n7274), .A3(n7273), .ZN(n7275) );
  NOR3_X1 U8522 ( .A1(n7276), .A2(n7275), .A3(n7280), .ZN(n7277) );
  OAI21_X1 U8523 ( .B1(n7278), .B2(n7277), .A(n7279), .ZN(n7284) );
  INV_X1 U8524 ( .A(n7279), .ZN(n7281) );
  OAI21_X1 U8525 ( .B1(n7281), .B2(n7280), .A(n7306), .ZN(n7283) );
  NOR3_X1 U8526 ( .A1(n9764), .A2(n7739), .A3(n9612), .ZN(n7282) );
  AOI21_X1 U8527 ( .B1(n7284), .B2(n7283), .A(n7282), .ZN(n7289) );
  INV_X1 U8528 ( .A(n7285), .ZN(n7287) );
  NOR2_X1 U8529 ( .A1(n9760), .A2(n9387), .ZN(n7286) );
  MUX2_X1 U8530 ( .A(n7287), .B(n7286), .S(n7739), .Z(n7288) );
  AOI21_X1 U8531 ( .B1(n7289), .B2(n9594), .A(n7288), .ZN(n7294) );
  NAND2_X1 U8532 ( .A1(n9589), .A2(n7306), .ZN(n7291) );
  NAND3_X1 U8533 ( .A1(n9756), .A2(n7739), .A3(n9386), .ZN(n7290) );
  OAI21_X1 U8534 ( .B1(n9756), .B2(n7291), .A(n7290), .ZN(n7293) );
  INV_X1 U8535 ( .A(n7292), .ZN(n7295) );
  OR2_X2 U8536 ( .A1(n7296), .A2(n7295), .ZN(n9566) );
  MUX2_X1 U8537 ( .A(n7296), .B(n7295), .S(n7739), .Z(n7297) );
  MUX2_X1 U8538 ( .A(n9748), .B(n10659), .S(n7739), .Z(n7300) );
  INV_X1 U8539 ( .A(n7300), .ZN(n7299) );
  MUX2_X1 U8540 ( .A(n9748), .B(n10659), .S(n7306), .Z(n7298) );
  NOR2_X1 U8541 ( .A1(n7301), .A2(n9260), .ZN(n7302) );
  NOR2_X1 U8542 ( .A1(n9744), .A2(n9384), .ZN(n7326) );
  NAND2_X1 U8543 ( .A1(n7303), .A2(n7739), .ZN(n7304) );
  AOI21_X1 U8544 ( .B1(n7322), .B2(n7304), .A(n7307), .ZN(n7305) );
  NAND2_X1 U8545 ( .A1(n7309), .A2(n7308), .ZN(n7311) );
  INV_X1 U8546 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9784) );
  OR2_X1 U8547 ( .A1(n6085), .A2(n9784), .ZN(n7310) );
  NAND2_X1 U8548 ( .A1(n7312), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7317) );
  INV_X1 U8549 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n7313) );
  OR2_X1 U8550 ( .A1(n6470), .A2(n7313), .ZN(n7316) );
  INV_X1 U8551 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7314) );
  OR2_X1 U8552 ( .A1(n5086), .A2(n7314), .ZN(n7315) );
  NAND4_X1 U8553 ( .A1(n7318), .A2(n7317), .A3(n7316), .A4(n7315), .ZN(n9535)
         );
  INV_X1 U8554 ( .A(n9535), .ZN(n7320) );
  AND2_X1 U8555 ( .A1(n9744), .A2(n9384), .ZN(n7349) );
  NOR2_X1 U8556 ( .A1(n7328), .A2(n7320), .ZN(n7327) );
  INV_X1 U8557 ( .A(n9744), .ZN(n7325) );
  AOI21_X1 U8558 ( .B1(n9741), .B2(n7325), .A(n7324), .ZN(n7329) );
  INV_X1 U8559 ( .A(n9594), .ZN(n7345) );
  XNOR2_X1 U8560 ( .A(n9764), .B(n9612), .ZN(n9604) );
  XNOR2_X1 U8561 ( .A(n9618), .B(n9601), .ZN(n9614) );
  INV_X1 U8562 ( .A(n8461), .ZN(n7340) );
  NOR4_X1 U8563 ( .A1(n5488), .A2(n7636), .A3(n8356), .A4(n7332), .ZN(n7333)
         );
  NAND4_X1 U8564 ( .A1(n7333), .A2(n7682), .A3(n7920), .A4(n7759), .ZN(n7334)
         );
  NOR4_X1 U8565 ( .A1(n7334), .A2(n6205), .A3(n7884), .A4(n8447), .ZN(n7338)
         );
  INV_X1 U8566 ( .A(n7335), .ZN(n7336) );
  OR2_X1 U8567 ( .A1(n7337), .A2(n7336), .ZN(n8322) );
  NAND4_X1 U8568 ( .A1(n6454), .A2(n8101), .A3(n7338), .A4(n8322), .ZN(n7339)
         );
  NOR4_X1 U8569 ( .A1(n8626), .A2(n8534), .A3(n7340), .A4(n7339), .ZN(n7341)
         );
  NAND3_X1 U8570 ( .A1(n8699), .A2(n8678), .A3(n7341), .ZN(n7342) );
  NOR4_X1 U8571 ( .A1(n5554), .A2(n8725), .A3(n6330), .A4(n7342), .ZN(n7343)
         );
  NAND4_X1 U8572 ( .A1(n9614), .A2(n9641), .A3(n7343), .A4(n9627), .ZN(n7344)
         );
  NOR4_X1 U8573 ( .A1(n9566), .A2(n7345), .A3(n9604), .A4(n7344), .ZN(n7346)
         );
  NAND3_X1 U8574 ( .A1(n7346), .A2(n9579), .A3(n9556), .ZN(n7347) );
  INV_X1 U8575 ( .A(n7350), .ZN(n7351) );
  OR2_X1 U8576 ( .A1(n7721), .A2(P2_U3151), .ZN(n8415) );
  INV_X1 U8577 ( .A(n7397), .ZN(n7352) );
  NOR3_X1 U8578 ( .A1(n7747), .A2(n7353), .A3(n5864), .ZN(n7356) );
  OAI21_X1 U8579 ( .B1(n8415), .B2(n7354), .A(P2_B_REG_SCAN_IN), .ZN(n7355) );
  OR2_X1 U8580 ( .A1(n7356), .A2(n7355), .ZN(n7357) );
  INV_X1 U8581 ( .A(n7358), .ZN(n7359) );
  INV_X2 U8582 ( .A(n10657), .ZN(P2_U3893) );
  NOR2_X1 U8583 ( .A1(n7362), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10582) );
  INV_X2 U8584 ( .A(n10582), .ZN(n8791) );
  OAI222_X1 U8585 ( .A1(n8793), .A2(n7360), .B1(n8791), .B2(n7364), .C1(
        P1_U3086), .C2(n7563), .ZN(P1_U3353) );
  NAND2_X1 U8586 ( .A1(n7361), .A2(P2_U3151), .ZN(n9261) );
  AND2_X1 U8587 ( .A1(n7362), .A2(P2_U3151), .ZN(n9787) );
  INV_X2 U8588 ( .A(n9787), .ZN(n9792) );
  OAI222_X1 U8589 ( .A1(n9261), .A2(n7365), .B1(n9792), .B2(n7364), .C1(
        P2_U3151), .C2(n7363), .ZN(P2_U3293) );
  INV_X1 U8590 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7367) );
  INV_X1 U8591 ( .A(n5868), .ZN(n7366) );
  OAI222_X1 U8592 ( .A1(n9261), .A2(n7367), .B1(n9792), .B2(n5115), .C1(
        P2_U3151), .C2(n7366), .ZN(P2_U3294) );
  OAI222_X1 U8593 ( .A1(n9261), .A2(n7368), .B1(n9792), .B2(n7384), .C1(
        P2_U3151), .C2(n7491), .ZN(P2_U3292) );
  OAI222_X1 U8594 ( .A1(n9261), .A2(n7370), .B1(n9792), .B2(n7378), .C1(
        P2_U3151), .C2(n7369), .ZN(P2_U3291) );
  OAI222_X1 U8595 ( .A1(n9261), .A2(n7372), .B1(n9792), .B2(n7381), .C1(
        P2_U3151), .C2(n7371), .ZN(P2_U3290) );
  OAI222_X1 U8596 ( .A1(n8793), .A2(n7373), .B1(n8791), .B2(n7375), .C1(
        P1_U3086), .C2(n7567), .ZN(P1_U3349) );
  OAI222_X1 U8597 ( .A1(n9261), .A2(n7376), .B1(n9792), .B2(n7375), .C1(
        P2_U3151), .C2(n7374), .ZN(P2_U3289) );
  OAI222_X1 U8598 ( .A1(n8793), .A2(n7377), .B1(n8791), .B2(n5115), .C1(
        P1_U3086), .C2(n7562), .ZN(P1_U3354) );
  OAI222_X1 U8599 ( .A1(n8793), .A2(n7379), .B1(n8791), .B2(n7378), .C1(
        P1_U3086), .C2(n7572), .ZN(P1_U3351) );
  OAI222_X1 U8600 ( .A1(n8793), .A2(n7382), .B1(n8791), .B2(n7381), .C1(
        P1_U3086), .C2(n7380), .ZN(P1_U3350) );
  OAI222_X1 U8601 ( .A1(n8793), .A2(n7385), .B1(n8791), .B2(n7384), .C1(
        P1_U3086), .C2(n7383), .ZN(P1_U3352) );
  INV_X1 U8602 ( .A(n9261), .ZN(n9790) );
  AOI22_X1 U8603 ( .A1(n10721), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n9790), .ZN(n7386) );
  OAI21_X1 U8604 ( .B1(n7388), .B2(n9792), .A(n7386), .ZN(P2_U3288) );
  OAI222_X1 U8605 ( .A1(n8793), .A2(n9187), .B1(n8791), .B2(n7388), .C1(
        P1_U3086), .C2(n7387), .ZN(P1_U3348) );
  INV_X1 U8606 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n7390) );
  NAND2_X1 U8607 ( .A1(n8238), .A2(n7397), .ZN(n7389) );
  OAI21_X1 U8608 ( .B1(n7397), .B2(n7390), .A(n7389), .ZN(P2_U3377) );
  INV_X1 U8609 ( .A(n7391), .ZN(n7395) );
  OAI222_X1 U8610 ( .A1(n9261), .A2(n7393), .B1(n9792), .B2(n7395), .C1(
        P2_U3151), .C2(n7392), .ZN(P2_U3287) );
  OAI222_X1 U8611 ( .A1(n8793), .A2(n7396), .B1(n8791), .B2(n7395), .C1(
        P1_U3086), .C2(n7394), .ZN(P1_U3347) );
  NAND2_X1 U8612 ( .A1(n6490), .A2(n7397), .ZN(n8786) );
  AND2_X1 U8613 ( .A1(n8786), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8614 ( .A1(n8786), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8615 ( .A1(n8786), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8616 ( .A1(n8786), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8617 ( .A1(n8786), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8618 ( .A1(n8786), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8619 ( .A1(n8786), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8620 ( .A1(n8786), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8621 ( .A1(n8786), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8622 ( .A1(n8786), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8623 ( .A1(n8786), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8624 ( .A1(n8786), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8625 ( .A1(n8786), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8626 ( .A1(n8786), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8627 ( .A1(n8786), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8628 ( .A1(n8786), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8629 ( .A1(n8786), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8630 ( .A1(n8786), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8631 ( .A1(n8786), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8632 ( .A1(n8786), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8633 ( .A1(n8786), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8634 ( .A1(n8786), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8635 ( .A1(n8786), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8636 ( .A1(n8786), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8637 ( .A1(n8786), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8638 ( .A1(n8786), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8639 ( .A1(n8786), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8640 ( .A1(n8786), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8641 ( .A1(n8786), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8642 ( .A1(n8786), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  INV_X1 U8643 ( .A(n7398), .ZN(n7402) );
  OAI222_X1 U8644 ( .A1(n9792), .A2(n7402), .B1(n8135), .B2(P2_U3151), .C1(
        n7399), .C2(n9783), .ZN(P2_U3286) );
  INV_X1 U8645 ( .A(n7400), .ZN(n7405) );
  INV_X1 U8646 ( .A(n8793), .ZN(n7822) );
  AOI22_X1 U8647 ( .A1(n10105), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n7822), .ZN(n7401) );
  OAI21_X1 U8648 ( .B1(n7405), .B2(n8791), .A(n7401), .ZN(P1_U3345) );
  INV_X1 U8649 ( .A(n8220), .ZN(n7881) );
  OAI222_X1 U8650 ( .A1(n8793), .A2(n9180), .B1(n8791), .B2(n7402), .C1(n7881), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8651 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7403) );
  OAI222_X1 U8652 ( .A1(n9792), .A2(n7405), .B1(n7404), .B2(P2_U3151), .C1(
        n7403), .C2(n9783), .ZN(P2_U3285) );
  MUX2_X1 U8653 ( .A(n9180), .B(n8449), .S(P2_U3893), .Z(n7406) );
  INV_X1 U8654 ( .A(n7406), .ZN(P2_U3500) );
  INV_X1 U8655 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7407) );
  OR2_X1 U8656 ( .A1(n8788), .A2(n10228), .ZN(n10750) );
  INV_X1 U8657 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n7574) );
  OAI22_X1 U8658 ( .A1(n7568), .A2(n7407), .B1(n10750), .B2(n7574), .ZN(n7408)
         );
  XNOR2_X1 U8659 ( .A(n7408), .B(P1_IR_REG_0__SCAN_IN), .ZN(n7415) );
  NAND2_X1 U8660 ( .A1(n7656), .A2(n7809), .ZN(n7409) );
  AND2_X1 U8661 ( .A1(n5090), .A2(n7409), .ZN(n7411) );
  INV_X1 U8662 ( .A(n7511), .ZN(n7519) );
  AOI21_X1 U8663 ( .B1(n7519), .B2(n7809), .A(P1_U3086), .ZN(n7412) );
  AND2_X1 U8664 ( .A1(n7411), .A2(n7412), .ZN(n7582) );
  INV_X1 U8665 ( .A(n7582), .ZN(n7569) );
  INV_X1 U8666 ( .A(n7411), .ZN(n7413) );
  AOI22_X1 U8667 ( .A1(n10756), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n7414) );
  OAI21_X1 U8668 ( .B1(n7415), .B2(n7569), .A(n7414), .ZN(P1_U3243) );
  INV_X1 U8669 ( .A(n7416), .ZN(n7419) );
  INV_X1 U8670 ( .A(n8390), .ZN(n7417) );
  OAI222_X1 U8671 ( .A1(n8793), .A2(n7418), .B1(n8791), .B2(n7419), .C1(
        P1_U3086), .C2(n7417), .ZN(P1_U3344) );
  OAI222_X1 U8672 ( .A1(n7420), .A2(P2_U3151), .B1(n9792), .B2(n7419), .C1(
        n9783), .C2(n5998), .ZN(P2_U3284) );
  NOR2_X1 U8673 ( .A1(n10756), .A2(P1_U3973), .ZN(P1_U3085) );
  MUX2_X1 U8674 ( .A(n7422), .B(n7421), .S(n5191), .Z(n7423) );
  NOR2_X1 U8675 ( .A1(n7423), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7424) );
  OAI22_X1 U8676 ( .A1(n7425), .A2(n10729), .B1(n10661), .B2(n7424), .ZN(n7426) );
  OAI21_X1 U8677 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n8357), .A(n7426), .ZN(n7427) );
  AOI21_X1 U8678 ( .B1(n9505), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n7427), .ZN(
        n7428) );
  OAI21_X1 U8679 ( .B1(n5904), .B2(n9521), .A(n7428), .ZN(P2_U3182) );
  NAND2_X1 U8680 ( .A1(n10104), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n7429) );
  OAI21_X1 U8681 ( .B1(n10433), .B2(n10104), .A(n7429), .ZN(P1_U3573) );
  INV_X1 U8682 ( .A(n7430), .ZN(n7434) );
  AOI22_X1 U8683 ( .A1(n8594), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n7822), .ZN(n7431) );
  OAI21_X1 U8684 ( .B1(n7434), .B2(n8791), .A(n7431), .ZN(P1_U3343) );
  INV_X1 U8685 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7432) );
  OAI222_X1 U8686 ( .A1(n9792), .A2(n7434), .B1(n7433), .B2(P2_U3151), .C1(
        n7432), .C2(n9783), .ZN(P2_U3283) );
  INV_X1 U8687 ( .A(n8746), .ZN(n8609) );
  NAND2_X1 U8688 ( .A1(n8609), .A2(P1_U3973), .ZN(n7435) );
  OAI21_X1 U8689 ( .B1(n5998), .B2(P1_U3973), .A(n7435), .ZN(P1_U3565) );
  INV_X1 U8690 ( .A(n10729), .ZN(n7453) );
  XNOR2_X1 U8691 ( .A(n7437), .B(n7436), .ZN(n7452) );
  INV_X1 U8692 ( .A(n9521), .ZN(n10722) );
  AOI21_X1 U8693 ( .B1(n7440), .B2(n7439), .A(n7438), .ZN(n7448) );
  AOI21_X1 U8694 ( .B1(n7443), .B2(n7442), .A(n7441), .ZN(n7444) );
  OAI22_X1 U8695 ( .A1(n10724), .A2(n7444), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8488), .ZN(n7445) );
  INV_X1 U8696 ( .A(n7445), .ZN(n7447) );
  NAND2_X1 U8697 ( .A1(n9505), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n7446) );
  OAI211_X1 U8698 ( .C1(n7448), .C2(n10717), .A(n7447), .B(n7446), .ZN(n7449)
         );
  AOI21_X1 U8699 ( .B1(n7450), .B2(n10722), .A(n7449), .ZN(n7451) );
  OAI21_X1 U8700 ( .B1(n7453), .B2(n7452), .A(n7451), .ZN(P2_U3184) );
  AOI21_X1 U8701 ( .B1(n7456), .B2(n7455), .A(n7454), .ZN(n7470) );
  XNOR2_X1 U8702 ( .A(n7458), .B(n7457), .ZN(n7459) );
  NAND2_X1 U8703 ( .A1(n7459), .A2(n10729), .ZN(n7469) );
  INV_X1 U8704 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7460) );
  NAND2_X1 U8705 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7786) );
  OAI21_X1 U8706 ( .B1(n10734), .B2(n7460), .A(n7786), .ZN(n7466) );
  AOI21_X1 U8707 ( .B1(n7463), .B2(n7462), .A(n7461), .ZN(n7464) );
  NOR2_X1 U8708 ( .A1(n7464), .A2(n10724), .ZN(n7465) );
  AOI211_X1 U8709 ( .C1(n10722), .C2(n7467), .A(n7466), .B(n7465), .ZN(n7468)
         );
  OAI211_X1 U8710 ( .C1(n7470), .C2(n10717), .A(n7469), .B(n7468), .ZN(
        P2_U3188) );
  INV_X1 U8711 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8966) );
  INV_X1 U8712 ( .A(n7471), .ZN(n7473) );
  OAI222_X1 U8713 ( .A1(n8793), .A2(n8966), .B1(n8791), .B2(n7473), .C1(
        P1_U3086), .C2(n10129), .ZN(P1_U3342) );
  INV_X1 U8714 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7474) );
  OAI222_X1 U8715 ( .A1(n9783), .A2(n7474), .B1(n9792), .B2(n7473), .C1(
        P2_U3151), .C2(n7472), .ZN(P2_U3282) );
  XNOR2_X1 U8716 ( .A(n7476), .B(n7475), .ZN(n7477) );
  NAND2_X1 U8717 ( .A1(n7477), .A2(n10729), .ZN(n7490) );
  AOI21_X1 U8718 ( .B1(n7480), .B2(n7479), .A(n7478), .ZN(n7481) );
  NOR2_X1 U8719 ( .A1(n10717), .A2(n7481), .ZN(n7488) );
  AOI21_X1 U8720 ( .B1(n8400), .B2(n7483), .A(n7482), .ZN(n7486) );
  INV_X1 U8721 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7484) );
  NOR2_X1 U8722 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7484), .ZN(n7753) );
  INV_X1 U8723 ( .A(n7753), .ZN(n7485) );
  OAI21_X1 U8724 ( .B1(n10724), .B2(n7486), .A(n7485), .ZN(n7487) );
  AOI211_X1 U8725 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n9505), .A(n7488), .B(
        n7487), .ZN(n7489) );
  OAI211_X1 U8726 ( .C1(n9521), .C2(n7491), .A(n7490), .B(n7489), .ZN(P2_U3185) );
  NAND2_X1 U8727 ( .A1(n8653), .A2(P1_B_REG_SCAN_IN), .ZN(n7493) );
  MUX2_X1 U8728 ( .A(n7493), .B(P1_B_REG_SCAN_IN), .S(n7492), .Z(n7494) );
  NAND2_X1 U8729 ( .A1(n8780), .A2(n8653), .ZN(n10575) );
  OAI21_X1 U8730 ( .B1(n10574), .B2(P1_D_REG_1__SCAN_IN), .A(n10575), .ZN(
        n7945) );
  NOR4_X1 U8731 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n7504) );
  NOR4_X1 U8732 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n7503) );
  OR4_X1 U8733 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_31__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n7501) );
  NOR4_X1 U8734 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n7499) );
  NOR4_X1 U8735 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n7498) );
  NOR4_X1 U8736 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n7497) );
  NOR4_X1 U8737 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n7496) );
  NAND4_X1 U8738 ( .A1(n7499), .A2(n7498), .A3(n7497), .A4(n7496), .ZN(n7500)
         );
  NOR4_X1 U8739 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n7501), .A4(n7500), .ZN(n7502) );
  AND3_X1 U8740 ( .A1(n7504), .A2(n7503), .A3(n7502), .ZN(n7505) );
  NOR2_X1 U8741 ( .A1(n10574), .A2(n7505), .ZN(n7536) );
  NOR2_X1 U8742 ( .A1(n7945), .A2(n7536), .ZN(n7506) );
  NAND2_X1 U8743 ( .A1(n8780), .A2(n8587), .ZN(n10576) );
  INV_X1 U8744 ( .A(n7946), .ZN(n7539) );
  AND2_X1 U8745 ( .A1(n7506), .A2(n7539), .ZN(n7528) );
  NAND2_X1 U8746 ( .A1(n7524), .A2(n5453), .ZN(n10041) );
  INV_X1 U8747 ( .A(n10087), .ZN(n10061) );
  INV_X1 U8748 ( .A(n7512), .ZN(n7513) );
  NAND2_X1 U8749 ( .A1(n7973), .A2(n9863), .ZN(n7514) );
  NAND2_X1 U8750 ( .A1(n7515), .A2(n7514), .ZN(n7644) );
  NAND2_X1 U8751 ( .A1(n7976), .A2(n9863), .ZN(n7516) );
  AOI21_X1 U8752 ( .B1(n5427), .B2(n7574), .A(n7511), .ZN(n7517) );
  NOR3_X1 U8753 ( .A1(n7644), .A2(n7518), .A3(n7517), .ZN(n7522) );
  NAND2_X1 U8754 ( .A1(n7518), .A2(n7644), .ZN(n7521) );
  NAND3_X1 U8755 ( .A1(n7519), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG1_REG_0__SCAN_IN), .ZN(n7520) );
  NAND2_X1 U8756 ( .A1(n7521), .A2(n7520), .ZN(n7646) );
  NOR2_X1 U8757 ( .A1(n7522), .A2(n7646), .ZN(n10751) );
  INV_X1 U8758 ( .A(n7161), .ZN(n8123) );
  NOR2_X1 U8759 ( .A1(n10557), .A2(n7656), .ZN(n7523) );
  NAND2_X1 U8760 ( .A1(n10751), .A2(n10081), .ZN(n7533) );
  AND2_X1 U8761 ( .A1(n7540), .A2(n7546), .ZN(n7951) );
  NAND2_X1 U8762 ( .A1(n7524), .A2(n7951), .ZN(n7527) );
  NAND2_X1 U8763 ( .A1(n10949), .A2(n7950), .ZN(n7537) );
  INV_X1 U8764 ( .A(n7537), .ZN(n7526) );
  INV_X1 U8765 ( .A(n7528), .ZN(n7531) );
  NAND2_X1 U8766 ( .A1(n7546), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8082) );
  NAND2_X1 U8767 ( .A1(n10557), .A2(n8082), .ZN(n7530) );
  NAND2_X1 U8768 ( .A1(n7656), .A2(n7508), .ZN(n7534) );
  INV_X1 U8769 ( .A(n7534), .ZN(n7529) );
  AOI21_X1 U8770 ( .B1(n7531), .B2(n7530), .A(n7529), .ZN(n7810) );
  NAND2_X1 U8771 ( .A1(n7810), .A2(n10573), .ZN(n8800) );
  AOI22_X1 U8772 ( .A1(n10073), .A2(n7976), .B1(n8800), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n7532) );
  OAI211_X1 U8773 ( .C1(n8799), .C2(n10061), .A(n7533), .B(n7532), .ZN(
        P1_U3232) );
  NAND2_X1 U8774 ( .A1(n10573), .A2(n7534), .ZN(n7535) );
  AND2_X1 U8775 ( .A1(n7945), .A2(n7537), .ZN(n7538) );
  INV_X1 U8776 ( .A(n7540), .ZN(n7550) );
  NAND2_X1 U8777 ( .A1(n7508), .A2(n7544), .ZN(n7545) );
  NAND2_X1 U8778 ( .A1(n7944), .A2(n7545), .ZN(n10848) );
  OR2_X1 U8779 ( .A1(n7547), .A2(n7546), .ZN(n10928) );
  OAI21_X1 U8780 ( .B1(n10821), .B2(n11022), .A(n7943), .ZN(n7549) );
  NOR2_X1 U8781 ( .A1(n8799), .A2(n10462), .ZN(n7942) );
  INV_X1 U8782 ( .A(n7942), .ZN(n7548) );
  OAI211_X1 U8783 ( .C1(n7977), .C2(n7550), .A(n7549), .B(n7548), .ZN(n7553)
         );
  NAND2_X1 U8784 ( .A1(n7553), .A2(n11037), .ZN(n7551) );
  OAI21_X1 U8785 ( .B1(n11037), .B2(n7574), .A(n7551), .ZN(P1_U3522) );
  INV_X1 U8786 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7555) );
  NAND2_X1 U8787 ( .A1(n7553), .A2(n11041), .ZN(n7554) );
  OAI21_X1 U8788 ( .B1(n11041), .B2(n7555), .A(n7554), .ZN(P1_U3453) );
  INV_X1 U8789 ( .A(n7556), .ZN(n7558) );
  OAI222_X1 U8790 ( .A1(n9783), .A2(n7557), .B1(n9792), .B2(n7558), .C1(
        P2_U3151), .C2(n9449), .ZN(P2_U3281) );
  OAI222_X1 U8791 ( .A1(n8793), .A2(n7559), .B1(n8791), .B2(n7558), .C1(
        P1_U3086), .C2(n10131), .ZN(P1_U3341) );
  NAND2_X1 U8792 ( .A1(n10380), .A2(P1_U3973), .ZN(n7560) );
  OAI21_X1 U8793 ( .B1(P1_U3973), .B2(n8417), .A(n7560), .ZN(P1_U3577) );
  INV_X1 U8794 ( .A(n7572), .ZN(n10769) );
  MUX2_X1 U8795 ( .A(n5425), .B(P1_REG2_REG_4__SCAN_IN), .S(n7572), .Z(n7561)
         );
  INV_X1 U8796 ( .A(n7561), .ZN(n10765) );
  NAND2_X1 U8797 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10650) );
  INV_X1 U8798 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7979) );
  AOI22_X1 U8799 ( .A1(n10654), .A2(n7979), .B1(P1_REG2_REG_1__SCAN_IN), .B2(
        n7562), .ZN(n10651) );
  NOR2_X1 U8800 ( .A1(n10650), .A2(n10651), .ZN(n10649) );
  AOI21_X1 U8801 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n10654), .A(n10649), .ZN(
        n10742) );
  INV_X1 U8802 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7564) );
  AOI22_X1 U8803 ( .A1(n10745), .A2(n7564), .B1(P1_REG2_REG_2__SCAN_IN), .B2(
        n7563), .ZN(n10741) );
  NOR2_X1 U8804 ( .A1(n10742), .A2(n10741), .ZN(n10740) );
  AOI21_X1 U8805 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n10745), .A(n10740), .ZN(
        n7590) );
  NAND2_X1 U8806 ( .A1(n7595), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7565) );
  OAI21_X1 U8807 ( .B1(n7595), .B2(P1_REG2_REG_3__SCAN_IN), .A(n7565), .ZN(
        n7591) );
  NOR2_X1 U8808 ( .A1(n7590), .A2(n7591), .ZN(n7589) );
  NAND2_X1 U8809 ( .A1(n7608), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7566) );
  OAI21_X1 U8810 ( .B1(n7608), .B2(P1_REG2_REG_5__SCAN_IN), .A(n7566), .ZN(
        n7603) );
  AOI21_X1 U8811 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n7608), .A(n7602), .ZN(
        n7571) );
  INV_X1 U8812 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n8005) );
  AOI22_X1 U8813 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(n7567), .B1(n7620), .B2(
        n8005), .ZN(n7570) );
  NOR2_X1 U8814 ( .A1(n7571), .A2(n7570), .ZN(n7615) );
  AOI211_X1 U8815 ( .C1(n7571), .C2(n7570), .A(n7615), .B(n10763), .ZN(n7588)
         );
  INV_X1 U8816 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10825) );
  MUX2_X1 U8817 ( .A(n10825), .B(P1_REG1_REG_4__SCAN_IN), .S(n7572), .Z(n10758) );
  NAND2_X1 U8818 ( .A1(n7595), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7577) );
  INV_X1 U8819 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7573) );
  MUX2_X1 U8820 ( .A(n7573), .B(P1_REG1_REG_1__SCAN_IN), .S(n10654), .Z(n10647) );
  NOR3_X1 U8821 ( .A1(n5427), .A2(n7574), .A3(n10647), .ZN(n10646) );
  AOI21_X1 U8822 ( .B1(n10654), .B2(P1_REG1_REG_1__SCAN_IN), .A(n10646), .ZN(
        n10739) );
  INV_X1 U8823 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7575) );
  MUX2_X1 U8824 ( .A(n7575), .B(P1_REG1_REG_2__SCAN_IN), .S(n10745), .Z(n10738) );
  NOR2_X1 U8825 ( .A1(n10739), .A2(n10738), .ZN(n10737) );
  AOI21_X1 U8826 ( .B1(n10745), .B2(P1_REG1_REG_2__SCAN_IN), .A(n10737), .ZN(
        n7594) );
  OAI21_X1 U8827 ( .B1(n7595), .B2(P1_REG1_REG_3__SCAN_IN), .A(n7577), .ZN(
        n7593) );
  NOR2_X1 U8828 ( .A1(n7594), .A2(n7593), .ZN(n7592) );
  INV_X1 U8829 ( .A(n7592), .ZN(n7576) );
  NAND2_X1 U8830 ( .A1(n7577), .A2(n7576), .ZN(n10757) );
  AND2_X1 U8831 ( .A1(n10758), .A2(n10757), .ZN(n10760) );
  AOI21_X1 U8832 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n10769), .A(n10760), .ZN(
        n7607) );
  NAND2_X1 U8833 ( .A1(n7608), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7578) );
  OAI21_X1 U8834 ( .B1(n7608), .B2(P1_REG1_REG_5__SCAN_IN), .A(n7578), .ZN(
        n7606) );
  NOR2_X1 U8835 ( .A1(n7607), .A2(n7606), .ZN(n7605) );
  AOI21_X1 U8836 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n7608), .A(n7605), .ZN(
        n7581) );
  INV_X1 U8837 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7579) );
  MUX2_X1 U8838 ( .A(n7579), .B(P1_REG1_REG_6__SCAN_IN), .S(n7620), .Z(n7580)
         );
  NOR2_X1 U8839 ( .A1(n7581), .A2(n7580), .ZN(n7619) );
  NAND2_X1 U8840 ( .A1(n7582), .A2(n7151), .ZN(n10759) );
  AOI211_X1 U8841 ( .C1(n7581), .C2(n7580), .A(n7619), .B(n10759), .ZN(n7587)
         );
  INV_X1 U8842 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n7585) );
  NAND2_X1 U8843 ( .A1(n7582), .A2(n8788), .ZN(n10220) );
  INV_X1 U8844 ( .A(n10220), .ZN(n10770) );
  NAND2_X1 U8845 ( .A1(n10770), .A2(n7620), .ZN(n7584) );
  NAND2_X1 U8846 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n7583) );
  OAI211_X1 U8847 ( .C1(n7585), .C2(n10203), .A(n7584), .B(n7583), .ZN(n7586)
         );
  OR3_X1 U8848 ( .A1(n7588), .A2(n7587), .A3(n7586), .ZN(P1_U3249) );
  AOI211_X1 U8849 ( .C1(n7591), .C2(n7590), .A(n7589), .B(n10763), .ZN(n7601)
         );
  AOI211_X1 U8850 ( .C1(n7594), .C2(n7593), .A(n7592), .B(n10759), .ZN(n7600)
         );
  INV_X1 U8851 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7598) );
  NAND2_X1 U8852 ( .A1(n10770), .A2(n7595), .ZN(n7597) );
  NAND2_X1 U8853 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n7596) );
  OAI211_X1 U8854 ( .C1(n7598), .C2(n10203), .A(n7597), .B(n7596), .ZN(n7599)
         );
  OR3_X1 U8855 ( .A1(n7601), .A2(n7600), .A3(n7599), .ZN(P1_U3246) );
  AOI211_X1 U8856 ( .C1(n7604), .C2(n7603), .A(n7602), .B(n10763), .ZN(n7614)
         );
  AOI211_X1 U8857 ( .C1(n7607), .C2(n7606), .A(n7605), .B(n10759), .ZN(n7613)
         );
  INV_X1 U8858 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7611) );
  NAND2_X1 U8859 ( .A1(n10770), .A2(n7608), .ZN(n7610) );
  NAND2_X1 U8860 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n7609) );
  OAI211_X1 U8861 ( .C1(n7611), .C2(n10203), .A(n7610), .B(n7609), .ZN(n7612)
         );
  OR3_X1 U8862 ( .A1(n7614), .A2(n7613), .A3(n7612), .ZN(P1_U3248) );
  AOI21_X1 U8863 ( .B1(n7620), .B2(P1_REG2_REG_6__SCAN_IN), .A(n7615), .ZN(
        n7618) );
  NAND2_X1 U8864 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n7706), .ZN(n7616) );
  OAI21_X1 U8865 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n7706), .A(n7616), .ZN(
        n7617) );
  NOR2_X1 U8866 ( .A1(n7618), .A2(n7617), .ZN(n7701) );
  AOI211_X1 U8867 ( .C1(n7618), .C2(n7617), .A(n7701), .B(n10763), .ZN(n7629)
         );
  AOI21_X1 U8868 ( .B1(n7620), .B2(P1_REG1_REG_6__SCAN_IN), .A(n7619), .ZN(
        n7623) );
  NAND2_X1 U8869 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n7706), .ZN(n7621) );
  OAI21_X1 U8870 ( .B1(n7706), .B2(P1_REG1_REG_7__SCAN_IN), .A(n7621), .ZN(
        n7622) );
  NOR2_X1 U8871 ( .A1(n7623), .A2(n7622), .ZN(n7705) );
  AOI211_X1 U8872 ( .C1(n7623), .C2(n7622), .A(n7705), .B(n10759), .ZN(n7628)
         );
  INV_X1 U8873 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7626) );
  NAND2_X1 U8874 ( .A1(n10770), .A2(n7706), .ZN(n7625) );
  NAND2_X1 U8875 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n7624) );
  OAI211_X1 U8876 ( .C1(n7626), .C2(n10203), .A(n7625), .B(n7624), .ZN(n7627)
         );
  OR3_X1 U8877 ( .A1(n7629), .A2(n7628), .A3(n7627), .ZN(P1_U3250) );
  NAND2_X1 U8878 ( .A1(n9718), .A2(n9653), .ZN(n7631) );
  NOR2_X1 U8879 ( .A1(n5619), .A2(n9637), .ZN(n8360) );
  AOI21_X1 U8880 ( .B1(n8356), .B2(n7631), .A(n8360), .ZN(n7678) );
  MUX2_X1 U8881 ( .A(n7421), .B(n7678), .S(n9735), .Z(n7632) );
  OAI21_X1 U8882 ( .B1(n7889), .B2(n9738), .A(n7632), .ZN(P2_U3459) );
  XNOR2_X1 U8883 ( .A(n7634), .B(n7633), .ZN(n8487) );
  NOR2_X1 U8884 ( .A1(n7930), .A2(n8726), .ZN(n8491) );
  XNOR2_X1 U8885 ( .A(n7636), .B(n7635), .ZN(n7637) );
  NAND2_X1 U8886 ( .A1(n7637), .A2(n9664), .ZN(n7639) );
  AOI22_X1 U8887 ( .A1(n9667), .A2(n9404), .B1(n9402), .B2(n9668), .ZN(n7638)
         );
  NAND2_X1 U8888 ( .A1(n7639), .A2(n7638), .ZN(n8489) );
  AOI211_X1 U8889 ( .C1(n8487), .C2(n9733), .A(n8491), .B(n8489), .ZN(n10802)
         );
  OR2_X1 U8890 ( .A1(n10802), .A2(n9683), .ZN(n7640) );
  OAI21_X1 U8891 ( .B1(n9735), .B2(n7641), .A(n7640), .ZN(P2_U3461) );
  INV_X1 U8892 ( .A(n7642), .ZN(n7663) );
  AOI22_X1 U8893 ( .A1(n10158), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n7822), .ZN(n7643) );
  OAI21_X1 U8894 ( .B1(n7663), .B2(n8791), .A(n7643), .ZN(P1_U3340) );
  NOR2_X1 U8895 ( .A1(n7644), .A2(n9951), .ZN(n7645) );
  NAND2_X1 U8896 ( .A1(n7077), .A2(n9863), .ZN(n7648) );
  NAND2_X1 U8897 ( .A1(n7649), .A2(n7648), .ZN(n7650) );
  XNOR2_X1 U8898 ( .A(n7650), .B(n9899), .ZN(n7651) );
  NAND2_X1 U8899 ( .A1(n7652), .A2(n7651), .ZN(n7795) );
  INV_X1 U8900 ( .A(n7651), .ZN(n7654) );
  INV_X1 U8901 ( .A(n7652), .ZN(n7653) );
  NAND2_X1 U8902 ( .A1(n7654), .A2(n7653), .ZN(n7794) );
  NAND2_X1 U8903 ( .A1(n7795), .A2(n7794), .ZN(n7655) );
  AOI22_X1 U8904 ( .A1(n7077), .A2(n9953), .B1(n7981), .B2(n9863), .ZN(n7793)
         );
  XNOR2_X1 U8905 ( .A(n7655), .B(n7793), .ZN(n7661) );
  INV_X1 U8906 ( .A(n7973), .ZN(n7658) );
  OAI22_X1 U8907 ( .A1(n7658), .A2(n10464), .B1(n7657), .B2(n10462), .ZN(n7971) );
  AOI22_X1 U8908 ( .A1(n7971), .A2(n10029), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n8800), .ZN(n7660) );
  NAND2_X1 U8909 ( .A1(n10073), .A2(n7981), .ZN(n7659) );
  OAI211_X1 U8910 ( .C1(n7661), .C2(n10064), .A(n7660), .B(n7659), .ZN(
        P1_U3222) );
  INV_X1 U8911 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7662) );
  OAI222_X1 U8912 ( .A1(n9792), .A2(n7663), .B1(n9466), .B2(P2_U3151), .C1(
        n7662), .C2(n9783), .ZN(P2_U3280) );
  OAI21_X1 U8913 ( .B1(n7665), .B2(n7667), .A(n7664), .ZN(n8404) );
  INV_X1 U8914 ( .A(n9401), .ZN(n8058) );
  INV_X1 U8915 ( .A(n9403), .ZN(n7751) );
  XNOR2_X1 U8916 ( .A(n7666), .B(n7667), .ZN(n7668) );
  OAI222_X1 U8917 ( .A1(n9637), .A2(n8058), .B1(n9635), .B2(n7751), .C1(n9653), 
        .C2(n7668), .ZN(n8399) );
  AOI21_X1 U8918 ( .B1(n9733), .B2(n8404), .A(n8399), .ZN(n7696) );
  INV_X1 U8919 ( .A(n9738), .ZN(n8453) );
  AOI22_X1 U8920 ( .A1(n8453), .A2(n7754), .B1(n9683), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n7669) );
  OAI21_X1 U8921 ( .B1(n7696), .B2(n9683), .A(n7669), .ZN(P2_U3462) );
  NAND2_X1 U8922 ( .A1(n7332), .A2(n7736), .ZN(n7670) );
  NAND2_X1 U8923 ( .A1(n7671), .A2(n7670), .ZN(n8249) );
  INV_X1 U8924 ( .A(n7672), .ZN(n7673) );
  XNOR2_X1 U8925 ( .A(n7332), .B(n7673), .ZN(n7676) );
  NAND2_X1 U8926 ( .A1(n8249), .A2(n8292), .ZN(n7675) );
  AOI22_X1 U8927 ( .A1(n9667), .A2(n9405), .B1(n9403), .B2(n9668), .ZN(n7674)
         );
  OAI211_X1 U8928 ( .C1(n9653), .C2(n7676), .A(n7675), .B(n7674), .ZN(n8246)
         );
  AOI21_X1 U8929 ( .B1(n6482), .B2(n8249), .A(n8246), .ZN(n7693) );
  AOI22_X1 U8930 ( .A1(n8453), .A2(n7733), .B1(n9683), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n7677) );
  OAI21_X1 U8931 ( .B1(n7693), .B2(n9683), .A(n7677), .ZN(P2_U3460) );
  MUX2_X1 U8932 ( .A(n6090), .B(n7678), .S(n11017), .Z(n7679) );
  OAI21_X1 U8933 ( .B1(n9779), .B2(n7889), .A(n7679), .ZN(P2_U3390) );
  OAI21_X1 U8934 ( .B1(n7681), .B2(n7682), .A(n7680), .ZN(n8316) );
  NOR2_X1 U8935 ( .A1(n8312), .A2(n8726), .ZN(n7687) );
  XNOR2_X1 U8936 ( .A(n7683), .B(n7682), .ZN(n7684) );
  NAND2_X1 U8937 ( .A1(n7684), .A2(n9664), .ZN(n7686) );
  AOI22_X1 U8938 ( .A1(n9668), .A2(n9400), .B1(n9402), .B2(n9667), .ZN(n7685)
         );
  NAND2_X1 U8939 ( .A1(n7686), .A2(n7685), .ZN(n8313) );
  AOI211_X1 U8940 ( .C1(n9733), .C2(n8316), .A(n7687), .B(n8313), .ZN(n10811)
         );
  OR2_X1 U8941 ( .A1(n10811), .A2(n9683), .ZN(n7688) );
  OAI21_X1 U8942 ( .B1(n9735), .B2(n6131), .A(n7688), .ZN(P2_U3463) );
  INV_X1 U8943 ( .A(n7689), .ZN(n7699) );
  AOI22_X1 U8944 ( .A1(n10182), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n7822), .ZN(n7690) );
  OAI21_X1 U8945 ( .B1(n7699), .B2(n8791), .A(n7690), .ZN(P1_U3339) );
  OAI22_X1 U8946 ( .A1(n9779), .A2(n8245), .B1(n11017), .B2(n6078), .ZN(n7691)
         );
  INV_X1 U8947 ( .A(n7691), .ZN(n7692) );
  OAI21_X1 U8948 ( .B1(n7693), .B2(n11015), .A(n7692), .ZN(P2_U3393) );
  OAI22_X1 U8949 ( .A1(n9779), .A2(n8401), .B1(n11017), .B2(n6117), .ZN(n7694)
         );
  INV_X1 U8950 ( .A(n7694), .ZN(n7695) );
  OAI21_X1 U8951 ( .B1(n7696), .B2(n11015), .A(n7695), .ZN(P2_U3399) );
  NAND2_X1 U8952 ( .A1(n10104), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7697) );
  OAI21_X1 U8953 ( .B1(n9960), .B2(n10104), .A(n7697), .ZN(P1_U3583) );
  OAI222_X1 U8954 ( .A1(n9261), .A2(n7700), .B1(n9792), .B2(n7699), .C1(
        P2_U3151), .C2(n7698), .ZN(P2_U3279) );
  NAND2_X1 U8955 ( .A1(n7873), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7702) );
  OAI21_X1 U8956 ( .B1(n7873), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7702), .ZN(
        n7703) );
  AOI211_X1 U8957 ( .C1(n7704), .C2(n7703), .A(n7872), .B(n10763), .ZN(n7715)
         );
  AOI21_X1 U8958 ( .B1(n7706), .B2(P1_REG1_REG_7__SCAN_IN), .A(n7705), .ZN(
        n7709) );
  NAND2_X1 U8959 ( .A1(n7873), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7707) );
  OAI21_X1 U8960 ( .B1(n7873), .B2(P1_REG1_REG_8__SCAN_IN), .A(n7707), .ZN(
        n7708) );
  NOR2_X1 U8961 ( .A1(n7709), .A2(n7708), .ZN(n7868) );
  AOI211_X1 U8962 ( .C1(n7709), .C2(n7708), .A(n7868), .B(n10759), .ZN(n7714)
         );
  INV_X1 U8963 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7712) );
  NAND2_X1 U8964 ( .A1(n10770), .A2(n7873), .ZN(n7711) );
  NAND2_X1 U8965 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n7710) );
  OAI211_X1 U8966 ( .C1(n7712), .C2(n10203), .A(n7711), .B(n7710), .ZN(n7713)
         );
  OR3_X1 U8967 ( .A1(n7715), .A2(n7714), .A3(n7713), .ZN(P1_U3251) );
  INV_X1 U8968 ( .A(n10305), .ZN(n9913) );
  NAND2_X1 U8969 ( .A1(n9913), .A2(P1_U3973), .ZN(n7716) );
  OAI21_X1 U8970 ( .B1(n6061), .B2(P1_U3973), .A(n7716), .ZN(P1_U3580) );
  INV_X1 U8971 ( .A(n7748), .ZN(n7728) );
  INV_X1 U8972 ( .A(n7717), .ZN(n7718) );
  NAND2_X1 U8973 ( .A1(n7746), .A2(n7718), .ZN(n7724) );
  INV_X1 U8974 ( .A(n7719), .ZN(n7720) );
  NAND2_X1 U8975 ( .A1(n7748), .A2(n7720), .ZN(n7723) );
  NAND4_X1 U8976 ( .A1(n7724), .A2(n7723), .A3(n7722), .A4(n7721), .ZN(n7738)
         );
  INV_X1 U8977 ( .A(n7725), .ZN(n7726) );
  OAI21_X1 U8978 ( .B1(n7738), .B2(n7726), .A(P2_STATE_REG_SCAN_IN), .ZN(n7727) );
  OAI21_X2 U8979 ( .B1(n7728), .B2(n7747), .A(n7727), .ZN(n9364) );
  OR2_X1 U8980 ( .A1(n7730), .A2(n7729), .ZN(n7732) );
  XNOR2_X1 U8981 ( .A(n7735), .B(n7733), .ZN(n7734) );
  OAI21_X1 U8982 ( .B1(n8363), .B2(n7766), .A(n7736), .ZN(n7935) );
  XNOR2_X1 U8983 ( .A(n7737), .B(n9403), .ZN(n7928) );
  NAND2_X1 U8984 ( .A1(n7927), .A2(n7928), .ZN(n7742) );
  NAND2_X1 U8985 ( .A1(n7737), .A2(n7751), .ZN(n7741) );
  AND2_X1 U8986 ( .A1(n7742), .A2(n7741), .ZN(n7744) );
  XNOR2_X1 U8987 ( .A(n7735), .B(n7754), .ZN(n7764) );
  XNOR2_X1 U8988 ( .A(n7764), .B(n7770), .ZN(n7743) );
  INV_X1 U8989 ( .A(n7738), .ZN(n7740) );
  OAI211_X1 U8990 ( .C1(n7744), .C2(n7743), .A(n5658), .B(n7765), .ZN(n7756)
         );
  OR2_X2 U8991 ( .A1(n7745), .A2(n7729), .ZN(n9590) );
  OAI21_X2 U8992 ( .B1(n7746), .B2(n7745), .A(n9590), .ZN(n9353) );
  INV_X1 U8993 ( .A(n9361), .ZN(n7750) );
  OAI22_X1 U8994 ( .A1(n9376), .A2(n7751), .B1(n8058), .B2(n9328), .ZN(n7752)
         );
  AOI211_X1 U8995 ( .C1(n7754), .C2(n9353), .A(n7753), .B(n7752), .ZN(n7755)
         );
  OAI211_X1 U8996 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n9377), .A(n7756), .B(
        n7755), .ZN(P2_U3158) );
  OAI21_X1 U8997 ( .B1(n7758), .B2(n7759), .A(n7757), .ZN(n8353) );
  NOR2_X1 U8998 ( .A1(n8349), .A2(n8726), .ZN(n7762) );
  INV_X1 U8999 ( .A(n9399), .ZN(n7964) );
  XNOR2_X1 U9000 ( .A(n7760), .B(n7759), .ZN(n7761) );
  OAI222_X1 U9001 ( .A1(n9637), .A2(n7964), .B1(n9635), .B2(n8058), .C1(n9653), 
        .C2(n7761), .ZN(n8350) );
  AOI211_X1 U9002 ( .C1(n9733), .C2(n8353), .A(n7762), .B(n8350), .ZN(n10836)
         );
  NAND2_X1 U9003 ( .A1(n9683), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7763) );
  OAI21_X1 U9004 ( .B1(n10836), .B2(n9683), .A(n7763), .ZN(P2_U3464) );
  AOI21_X1 U9005 ( .B1(n7768), .B2(n7767), .A(n7778), .ZN(n7776) );
  INV_X1 U9006 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7769) );
  NOR2_X1 U9007 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7769), .ZN(n10681) );
  INV_X1 U9008 ( .A(n9400), .ZN(n7922) );
  OAI22_X1 U9009 ( .A1(n9376), .A2(n7770), .B1(n7922), .B2(n9328), .ZN(n7771)
         );
  AOI211_X1 U9010 ( .C1(n7772), .C2(n9353), .A(n10681), .B(n7771), .ZN(n7775)
         );
  INV_X1 U9011 ( .A(n8311), .ZN(n7773) );
  NAND2_X1 U9012 ( .A1(n9364), .A2(n7773), .ZN(n7774) );
  OAI211_X1 U9013 ( .C1(n7776), .C2(n9355), .A(n7775), .B(n7774), .ZN(P2_U3170) );
  XNOR2_X1 U9014 ( .A(n8831), .B(n7779), .ZN(n7780) );
  XNOR2_X1 U9015 ( .A(n7780), .B(n9400), .ZN(n8056) );
  NOR2_X1 U9016 ( .A1(n7780), .A2(n9400), .ZN(n7784) );
  INV_X1 U9017 ( .A(n7784), .ZN(n7782) );
  XNOR2_X1 U9018 ( .A(n7735), .B(n7790), .ZN(n7957) );
  XNOR2_X1 U9019 ( .A(n7957), .B(n9399), .ZN(n7783) );
  INV_X1 U9020 ( .A(n7783), .ZN(n7781) );
  OAI21_X1 U9021 ( .B1(n8055), .B2(n7784), .A(n7783), .ZN(n7785) );
  NAND3_X1 U9022 ( .A1(n5644), .A2(n5658), .A3(n7785), .ZN(n7792) );
  INV_X1 U9023 ( .A(n7786), .ZN(n7787) );
  AOI21_X1 U9024 ( .B1(n9380), .B2(n9398), .A(n7787), .ZN(n7788) );
  OAI21_X1 U9025 ( .B1(n7922), .B2(n9376), .A(n7788), .ZN(n7789) );
  AOI21_X1 U9026 ( .B1(n7790), .B2(n9353), .A(n7789), .ZN(n7791) );
  OAI211_X1 U9027 ( .C1(n8409), .C2(n9377), .A(n7792), .B(n7791), .ZN(P2_U3179) );
  NAND2_X1 U9028 ( .A1(n7794), .A2(n7793), .ZN(n7796) );
  NAND2_X1 U9029 ( .A1(n7796), .A2(n7795), .ZN(n8795) );
  OAI22_X1 U9030 ( .A1(n7799), .A2(n9860), .B1(n7657), .B2(n7808), .ZN(n7798)
         );
  XNOR2_X1 U9031 ( .A(n7798), .B(n9899), .ZN(n7802) );
  OR2_X1 U9032 ( .A1(n7657), .A2(n9901), .ZN(n7801) );
  INV_X1 U9033 ( .A(n7799), .ZN(n10795) );
  NAND2_X1 U9034 ( .A1(n10795), .A2(n9863), .ZN(n7800) );
  NAND2_X1 U9035 ( .A1(n7801), .A2(n7800), .ZN(n7803) );
  XNOR2_X1 U9036 ( .A(n7802), .B(n7803), .ZN(n8796) );
  INV_X1 U9037 ( .A(n7803), .ZN(n7804) );
  NAND2_X1 U9038 ( .A1(n7802), .A2(n7804), .ZN(n7805) );
  OAI22_X1 U9039 ( .A1(n8798), .A2(n7808), .B1(n7806), .B2(n9860), .ZN(n7807)
         );
  XNOR2_X1 U9040 ( .A(n7807), .B(n9899), .ZN(n7826) );
  OAI22_X1 U9041 ( .A1(n8798), .A2(n9901), .B1(n7806), .B2(n7808), .ZN(n7827)
         );
  XNOR2_X1 U9042 ( .A(n7826), .B(n7827), .ZN(n7824) );
  XNOR2_X1 U9043 ( .A(n7825), .B(n7824), .ZN(n7815) );
  NAND3_X1 U9044 ( .A1(n7810), .A2(n7511), .A3(n7809), .ZN(n7811) );
  MUX2_X1 U9045 ( .A(P1_U3086), .B(n10071), .S(n8033), .Z(n7814) );
  AOI22_X1 U9046 ( .A1(n10550), .A2(n7812), .B1(n10102), .B2(n10552), .ZN(
        n8029) );
  OAI22_X1 U9047 ( .A1(n8029), .A2(n10041), .B1(n7806), .B2(n10090), .ZN(n7813) );
  AOI211_X1 U9048 ( .C1(n7815), .C2(n10081), .A(n7814), .B(n7813), .ZN(n7816)
         );
  INV_X1 U9049 ( .A(n7816), .ZN(P1_U3218) );
  INV_X1 U9050 ( .A(n7817), .ZN(n7820) );
  AOI22_X1 U9051 ( .A1(n10198), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n7822), .ZN(n7818) );
  OAI21_X1 U9052 ( .B1(n7820), .B2(n8791), .A(n7818), .ZN(P1_U3338) );
  OAI222_X1 U9053 ( .A1(n9792), .A2(n7820), .B1(n9506), .B2(P2_U3151), .C1(
        n7819), .C2(n9783), .ZN(P2_U3278) );
  INV_X1 U9054 ( .A(n7821), .ZN(n7865) );
  AOI22_X1 U9055 ( .A1(n10209), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n7822), .ZN(n7823) );
  OAI21_X1 U9056 ( .B1(n7865), .B2(n8791), .A(n7823), .ZN(P1_U3337) );
  INV_X1 U9057 ( .A(n10828), .ZN(n7844) );
  INV_X1 U9058 ( .A(n7826), .ZN(n7828) );
  OR2_X1 U9059 ( .A1(n7828), .A2(n7827), .ZN(n7829) );
  OAI22_X1 U9060 ( .A1(n8015), .A2(n7808), .B1(n10816), .B2(n9860), .ZN(n7830)
         );
  XNOR2_X1 U9061 ( .A(n7830), .B(n9951), .ZN(n7833) );
  OR2_X1 U9062 ( .A1(n8015), .A2(n9901), .ZN(n7832) );
  INV_X2 U9063 ( .A(n7808), .ZN(n9954) );
  NAND2_X1 U9064 ( .A1(n10829), .A2(n9954), .ZN(n7831) );
  NAND2_X1 U9065 ( .A1(n7832), .A2(n7831), .ZN(n7834) );
  NAND2_X1 U9066 ( .A1(n7833), .A2(n7834), .ZN(n8064) );
  INV_X1 U9067 ( .A(n7833), .ZN(n7836) );
  INV_X1 U9068 ( .A(n7834), .ZN(n7835) );
  NAND2_X1 U9069 ( .A1(n7836), .A2(n7835), .ZN(n7837) );
  NAND2_X1 U9070 ( .A1(n8064), .A2(n7837), .ZN(n7839) );
  AOI21_X1 U9071 ( .B1(n7838), .B2(n7839), .A(n10064), .ZN(n7840) );
  NAND2_X1 U9072 ( .A1(n7840), .A2(n8065), .ZN(n7843) );
  AOI22_X1 U9073 ( .A1(n10550), .A2(n10103), .B1(n10101), .B2(n10552), .ZN(
        n10819) );
  NAND2_X1 U9074 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10754) );
  OAI21_X1 U9075 ( .B1(n10819), .B2(n10041), .A(n10754), .ZN(n7841) );
  AOI21_X1 U9076 ( .B1(n10829), .B2(n10073), .A(n7841), .ZN(n7842) );
  OAI211_X1 U9077 ( .C1(n10084), .C2(n7844), .A(n7843), .B(n7842), .ZN(
        P1_U3230) );
  AOI21_X1 U9078 ( .B1(n7847), .B2(n7846), .A(n7845), .ZN(n7864) );
  INV_X1 U9079 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7855) );
  NOR2_X1 U9080 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7848), .ZN(n8050) );
  INV_X1 U9081 ( .A(n8050), .ZN(n7854) );
  AND2_X1 U9082 ( .A1(n7850), .A2(n7849), .ZN(n7852) );
  OAI21_X1 U9083 ( .B1(n7852), .B2(n7851), .A(n10729), .ZN(n7853) );
  OAI211_X1 U9084 ( .C1(n10734), .C2(n7855), .A(n7854), .B(n7853), .ZN(n7861)
         );
  AOI21_X1 U9085 ( .B1(n7858), .B2(n7857), .A(n7856), .ZN(n7859) );
  NOR2_X1 U9086 ( .A1(n7859), .A2(n10717), .ZN(n7860) );
  AOI211_X1 U9087 ( .C1(n10722), .C2(n7862), .A(n7861), .B(n7860), .ZN(n7863)
         );
  OAI21_X1 U9088 ( .B1(n7864), .B2(n10724), .A(n7863), .ZN(P2_U3190) );
  INV_X1 U9089 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7866) );
  OAI222_X1 U9090 ( .A1(n9261), .A2(n7866), .B1(P2_U3151), .B2(n9522), .C1(
        n7865), .C2(n9792), .ZN(P2_U3277) );
  INV_X1 U9091 ( .A(n10759), .ZN(n10147) );
  NOR2_X1 U9092 ( .A1(n8220), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7867) );
  AOI21_X1 U9093 ( .B1(n8220), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7867), .ZN(
        n7870) );
  AOI21_X1 U9094 ( .B1(n7873), .B2(P1_REG1_REG_8__SCAN_IN), .A(n7868), .ZN(
        n7869) );
  NAND2_X1 U9095 ( .A1(n7870), .A2(n7869), .ZN(n8221) );
  OAI21_X1 U9096 ( .B1(n7870), .B2(n7869), .A(n8221), .ZN(n7877) );
  NOR2_X1 U9097 ( .A1(n8220), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7871) );
  AOI21_X1 U9098 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n8220), .A(n7871), .ZN(
        n7875) );
  OAI21_X1 U9099 ( .B1(n7875), .B2(n7874), .A(n8215), .ZN(n7876) );
  AOI22_X1 U9100 ( .A1(n10147), .A2(n7877), .B1(n10222), .B2(n7876), .ZN(n7880) );
  NAND2_X1 U9101 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n8341) );
  INV_X1 U9102 ( .A(n8341), .ZN(n7878) );
  AOI21_X1 U9103 ( .B1(n10756), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7878), .ZN(
        n7879) );
  OAI211_X1 U9104 ( .C1(n7881), .C2(n10220), .A(n7880), .B(n7879), .ZN(
        P1_U3252) );
  OAI21_X1 U9105 ( .B1(n7883), .B2(n6451), .A(n7882), .ZN(n10867) );
  XNOR2_X1 U9106 ( .A(n7885), .B(n7884), .ZN(n7886) );
  AOI222_X1 U9107 ( .A1(n9664), .A2(n7886), .B1(n9397), .B2(n9668), .C1(n9399), 
        .C2(n9667), .ZN(n10866) );
  OAI21_X1 U9108 ( .B1(n9718), .B2(n10867), .A(n10866), .ZN(n7913) );
  INV_X1 U9109 ( .A(n7913), .ZN(n7888) );
  AOI22_X1 U9110 ( .A1(n8453), .A2(n10870), .B1(n9683), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n7887) );
  OAI21_X1 U9111 ( .B1(n7888), .B2(n9683), .A(n7887), .ZN(P2_U3466) );
  NOR2_X1 U9112 ( .A1(n9364), .A2(P2_U3151), .ZN(n7941) );
  INV_X1 U9113 ( .A(n9353), .ZN(n9383) );
  OAI22_X1 U9114 ( .A1(n9383), .A2(n7889), .B1(n9328), .B2(n5619), .ZN(n7890)
         );
  AOI21_X1 U9115 ( .B1(n5658), .B2(n8356), .A(n7890), .ZN(n7891) );
  OAI21_X1 U9116 ( .B1(n7941), .B2(n8357), .A(n7891), .ZN(P2_U3172) );
  NOR2_X1 U9117 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n7892) );
  AOI21_X1 U9118 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n7892), .ZN(n10645) );
  NOR2_X1 U9119 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7893) );
  AOI21_X1 U9120 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7893), .ZN(n10642) );
  INV_X1 U9121 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10165) );
  INV_X1 U9122 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9487) );
  AOI22_X1 U9123 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .B1(n10165), .B2(n9487), .ZN(n10639) );
  NOR2_X1 U9124 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7894) );
  AOI21_X1 U9125 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7894), .ZN(n10636) );
  NOR2_X1 U9126 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7895) );
  AOI21_X1 U9127 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7895), .ZN(n10633) );
  NOR2_X1 U9128 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7896) );
  AOI21_X1 U9129 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7896), .ZN(n10630) );
  NOR2_X1 U9130 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7897) );
  AOI21_X1 U9131 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7897), .ZN(n10627) );
  NOR2_X1 U9132 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7898) );
  AOI21_X1 U9133 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7898), .ZN(n10624) );
  NOR2_X1 U9134 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7899) );
  AOI21_X1 U9135 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7899), .ZN(n10621) );
  NOR2_X1 U9136 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7900) );
  AOI21_X1 U9137 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7900), .ZN(n10618) );
  NOR2_X1 U9138 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7901) );
  AOI21_X1 U9139 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7901), .ZN(n10615) );
  NOR2_X1 U9140 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7902) );
  AOI21_X1 U9141 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7902), .ZN(n10612) );
  NOR2_X1 U9142 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7903) );
  AOI21_X1 U9143 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7903), .ZN(n10609) );
  NOR2_X1 U9144 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7904) );
  AOI21_X1 U9145 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7904), .ZN(n10606) );
  AND2_X1 U9146 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n7905) );
  NOR2_X1 U9147 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7905), .ZN(n10592) );
  INV_X1 U9148 ( .A(n10592), .ZN(n10593) );
  INV_X1 U9149 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10674) );
  NAND3_X1 U9150 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10594) );
  NAND2_X1 U9151 ( .A1(n10674), .A2(n10594), .ZN(n10591) );
  NAND2_X1 U9152 ( .A1(n10593), .A2(n10591), .ZN(n10597) );
  NAND2_X1 U9153 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7906) );
  OAI21_X1 U9154 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7906), .ZN(n10596) );
  NOR2_X1 U9155 ( .A1(n10597), .A2(n10596), .ZN(n10595) );
  AOI21_X1 U9156 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10595), .ZN(n10600) );
  NAND2_X1 U9157 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7907) );
  OAI21_X1 U9158 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n7907), .ZN(n10599) );
  NOR2_X1 U9159 ( .A1(n10600), .A2(n10599), .ZN(n10598) );
  AOI21_X1 U9160 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10598), .ZN(n10603) );
  NOR2_X1 U9161 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7908) );
  AOI21_X1 U9162 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7908), .ZN(n10602) );
  NAND2_X1 U9163 ( .A1(n10603), .A2(n10602), .ZN(n10601) );
  OAI21_X1 U9164 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10601), .ZN(n10605) );
  NAND2_X1 U9165 ( .A1(n10606), .A2(n10605), .ZN(n10604) );
  OAI21_X1 U9166 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10604), .ZN(n10608) );
  NAND2_X1 U9167 ( .A1(n10609), .A2(n10608), .ZN(n10607) );
  OAI21_X1 U9168 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10607), .ZN(n10611) );
  NAND2_X1 U9169 ( .A1(n10612), .A2(n10611), .ZN(n10610) );
  OAI21_X1 U9170 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10610), .ZN(n10614) );
  NAND2_X1 U9171 ( .A1(n10615), .A2(n10614), .ZN(n10613) );
  OAI21_X1 U9172 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10613), .ZN(n10617) );
  NAND2_X1 U9173 ( .A1(n10618), .A2(n10617), .ZN(n10616) );
  OAI21_X1 U9174 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10616), .ZN(n10620) );
  NAND2_X1 U9175 ( .A1(n10621), .A2(n10620), .ZN(n10619) );
  OAI21_X1 U9176 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10619), .ZN(n10623) );
  NAND2_X1 U9177 ( .A1(n10624), .A2(n10623), .ZN(n10622) );
  OAI21_X1 U9178 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10622), .ZN(n10626) );
  NAND2_X1 U9179 ( .A1(n10627), .A2(n10626), .ZN(n10625) );
  OAI21_X1 U9180 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10625), .ZN(n10629) );
  NAND2_X1 U9181 ( .A1(n10630), .A2(n10629), .ZN(n10628) );
  OAI21_X1 U9182 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10628), .ZN(n10632) );
  NAND2_X1 U9183 ( .A1(n10633), .A2(n10632), .ZN(n10631) );
  OAI21_X1 U9184 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10631), .ZN(n10635) );
  NAND2_X1 U9185 ( .A1(n10636), .A2(n10635), .ZN(n10634) );
  OAI21_X1 U9186 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10634), .ZN(n10638) );
  NAND2_X1 U9187 ( .A1(n10639), .A2(n10638), .ZN(n10637) );
  OAI21_X1 U9188 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10637), .ZN(n10641) );
  NAND2_X1 U9189 ( .A1(n10642), .A2(n10641), .ZN(n10640) );
  OAI21_X1 U9190 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10640), .ZN(n10644) );
  NAND2_X1 U9191 ( .A1(n10645), .A2(n10644), .ZN(n10643) );
  OAI21_X1 U9192 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10643), .ZN(n7911) );
  XNOR2_X1 U9193 ( .A(n7909), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7910) );
  XNOR2_X1 U9194 ( .A(n7911), .B(n7910), .ZN(ADD_1068_U4) );
  OAI22_X1 U9195 ( .A1(n9779), .A2(n7968), .B1(n11017), .B2(n6166), .ZN(n7912)
         );
  AOI21_X1 U9196 ( .B1(n7913), .B2(n11017), .A(n7912), .ZN(n7914) );
  INV_X1 U9197 ( .A(n7914), .ZN(P2_U3411) );
  INV_X1 U9198 ( .A(n7920), .ZN(n7916) );
  NAND3_X1 U9199 ( .A1(n7757), .A2(n7917), .A3(n7916), .ZN(n7918) );
  NAND2_X1 U9200 ( .A1(n7915), .A2(n7918), .ZN(n8412) );
  NOR2_X1 U9201 ( .A1(n8408), .A2(n8726), .ZN(n7923) );
  XOR2_X1 U9202 ( .A(n7920), .B(n7919), .Z(n7921) );
  OAI222_X1 U9203 ( .A1(n9637), .A2(n5647), .B1(n9635), .B2(n7922), .C1(n7921), 
        .C2(n9653), .ZN(n8407) );
  AOI211_X1 U9204 ( .C1(n9733), .C2(n8412), .A(n7923), .B(n8407), .ZN(n10846)
         );
  OR2_X1 U9205 ( .A1(n10846), .A2(n9683), .ZN(n7924) );
  OAI21_X1 U9206 ( .B1(n9735), .B2(n7925), .A(n7924), .ZN(P2_U3465) );
  NAND2_X1 U9207 ( .A1(n10657), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7926) );
  OAI21_X1 U9208 ( .B1(n9550), .B2(n10657), .A(n7926), .ZN(P2_U3520) );
  OAI21_X1 U9209 ( .B1(n7928), .B2(n7927), .A(n7742), .ZN(n7929) );
  NAND2_X1 U9210 ( .A1(n7929), .A2(n5658), .ZN(n7933) );
  OAI22_X1 U9211 ( .A1(n9376), .A2(n5619), .B1(n7930), .B2(n9383), .ZN(n7931)
         );
  AOI21_X1 U9212 ( .B1(n9380), .B2(n9402), .A(n7931), .ZN(n7932) );
  OAI211_X1 U9213 ( .C1(n7941), .C2(n8488), .A(n7933), .B(n7932), .ZN(P2_U3177) );
  OAI21_X1 U9214 ( .B1(n7936), .B2(n7935), .A(n7934), .ZN(n7937) );
  NAND2_X1 U9215 ( .A1(n7937), .A2(n5658), .ZN(n7940) );
  OAI22_X1 U9216 ( .A1(n9376), .A2(n6447), .B1(n9383), .B2(n8245), .ZN(n7938)
         );
  AOI21_X1 U9217 ( .B1(n9380), .B2(n9403), .A(n7938), .ZN(n7939) );
  OAI211_X1 U9218 ( .C1(n7941), .C2(n8244), .A(n7940), .B(n7939), .ZN(P2_U3162) );
  AOI21_X1 U9219 ( .B1(n7944), .B2(n7943), .A(n7942), .ZN(n7955) );
  INV_X1 U9220 ( .A(n7945), .ZN(n7947) );
  NAND3_X1 U9221 ( .A1(n7948), .A2(n7947), .A3(n7946), .ZN(n7949) );
  AOI22_X1 U9222 ( .A1(n10955), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n10992), .ZN(n7954) );
  NOR2_X2 U9223 ( .A1(n10955), .A2(n7950), .ZN(n10959) );
  INV_X1 U9224 ( .A(n10949), .ZN(n10976) );
  NOR2_X1 U9225 ( .A1(n10477), .A2(n10976), .ZN(n11001) );
  INV_X1 U9226 ( .A(n7951), .ZN(n7952) );
  OAI21_X1 U9227 ( .B1(n11001), .B2(n10956), .A(n7976), .ZN(n7953) );
  OAI211_X1 U9228 ( .C1(n7955), .C2(n10955), .A(n7954), .B(n7953), .ZN(
        P1_U3293) );
  INV_X1 U9229 ( .A(n7766), .ZN(n8831) );
  XNOR2_X1 U9230 ( .A(n7968), .B(n8831), .ZN(n8045) );
  XNOR2_X1 U9231 ( .A(n8045), .B(n9398), .ZN(n7959) );
  OAI21_X1 U9232 ( .B1(n7959), .B2(n7958), .A(n8046), .ZN(n7960) );
  NAND2_X1 U9233 ( .A1(n7960), .A2(n5658), .ZN(n7967) );
  INV_X1 U9234 ( .A(n7961), .ZN(n10872) );
  INV_X1 U9235 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7962) );
  NOR2_X1 U9236 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7962), .ZN(n10720) );
  AOI21_X1 U9237 ( .B1(n9380), .B2(n9397), .A(n10720), .ZN(n7963) );
  OAI21_X1 U9238 ( .B1(n7964), .B2(n9376), .A(n7963), .ZN(n7965) );
  AOI21_X1 U9239 ( .B1(n10872), .B2(n9364), .A(n7965), .ZN(n7966) );
  OAI211_X1 U9240 ( .C1(n7968), .C2(n9383), .A(n7967), .B(n7966), .ZN(P2_U3153) );
  XNOR2_X1 U9241 ( .A(n7969), .B(n7970), .ZN(n7972) );
  AOI21_X1 U9242 ( .B1(n7972), .B2(n10821), .A(n7971), .ZN(n10775) );
  NAND2_X1 U9243 ( .A1(n7973), .A2(n7976), .ZN(n7990) );
  XNOR2_X1 U9244 ( .A(n7990), .B(n7969), .ZN(n10777) );
  INV_X1 U9245 ( .A(n10777), .ZN(n7984) );
  NAND2_X1 U9246 ( .A1(n10475), .A2(n10990), .ZN(n7975) );
  OR2_X1 U9247 ( .A1(n11005), .A2(n7974), .ZN(n10997) );
  OR2_X1 U9248 ( .A1(n7981), .A2(n7976), .ZN(n10784) );
  OAI211_X1 U9249 ( .C1(n7977), .C2(n10776), .A(n10949), .B(n10784), .ZN(
        n10774) );
  INV_X1 U9250 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7978) );
  OAI22_X1 U9251 ( .A1(n10475), .A2(n7979), .B1(n7978), .B2(n10472), .ZN(n7980) );
  AOI21_X1 U9252 ( .B1(n10956), .B2(n7981), .A(n7980), .ZN(n7982) );
  OAI21_X1 U9253 ( .B1(n10477), .B2(n10774), .A(n7982), .ZN(n7983) );
  AOI21_X1 U9254 ( .B1(n7984), .B2(n10961), .A(n7983), .ZN(n7985) );
  OAI21_X1 U9255 ( .B1(n10775), .B2(n11005), .A(n7985), .ZN(P1_U3292) );
  NAND2_X1 U9256 ( .A1(n7987), .A2(n7986), .ZN(n8179) );
  XOR2_X1 U9257 ( .A(n8179), .B(n7988), .Z(n7989) );
  OAI22_X1 U9258 ( .A1(n5344), .A2(n10462), .B1(n8071), .B2(n10464), .ZN(n8163) );
  AOI21_X1 U9259 ( .B1(n7989), .B2(n10821), .A(n8163), .ZN(n10850) );
  NAND2_X1 U9260 ( .A1(n7991), .A2(n7990), .ZN(n7993) );
  NAND2_X1 U9261 ( .A1(n8799), .A2(n10776), .ZN(n7992) );
  NAND2_X1 U9262 ( .A1(n7993), .A2(n7992), .ZN(n10782) );
  NAND2_X1 U9263 ( .A1(n10782), .A2(n10783), .ZN(n7995) );
  NAND2_X1 U9264 ( .A1(n7657), .A2(n7799), .ZN(n7994) );
  NAND2_X1 U9265 ( .A1(n7995), .A2(n7994), .ZN(n8031) );
  NAND2_X1 U9266 ( .A1(n8031), .A2(n8032), .ZN(n7997) );
  NAND2_X1 U9267 ( .A1(n8798), .A2(n7806), .ZN(n7996) );
  NAND2_X1 U9268 ( .A1(n7997), .A2(n7996), .ZN(n10812) );
  NAND2_X1 U9269 ( .A1(n10812), .A2(n10818), .ZN(n7999) );
  NAND2_X1 U9270 ( .A1(n8015), .A2(n10816), .ZN(n7998) );
  NAND2_X1 U9271 ( .A1(n7999), .A2(n7998), .ZN(n8019) );
  NAND2_X1 U9272 ( .A1(n8019), .A2(n8020), .ZN(n8001) );
  NAND2_X1 U9273 ( .A1(n8071), .A2(n10838), .ZN(n8000) );
  NAND2_X1 U9274 ( .A1(n8001), .A2(n8000), .ZN(n8180) );
  XOR2_X1 U9275 ( .A(n8179), .B(n8180), .Z(n10847) );
  INV_X1 U9276 ( .A(n10847), .ZN(n8009) );
  INV_X1 U9277 ( .A(n8189), .ZN(n8003) );
  OAI211_X1 U9278 ( .C1(n8002), .C2(n8022), .A(n8003), .B(n10949), .ZN(n10849)
         );
  INV_X1 U9279 ( .A(n8166), .ZN(n8004) );
  OAI22_X1 U9280 ( .A1(n10475), .A2(n8005), .B1(n8004), .B2(n10472), .ZN(n8006) );
  AOI21_X1 U9281 ( .B1(n10956), .B2(n8149), .A(n8006), .ZN(n8007) );
  OAI21_X1 U9282 ( .B1(n10849), .B2(n10477), .A(n8007), .ZN(n8008) );
  AOI21_X1 U9283 ( .B1(n8009), .B2(n10961), .A(n8008), .ZN(n8010) );
  OAI21_X1 U9284 ( .B1(n10955), .B2(n10850), .A(n8010), .ZN(P1_U3287) );
  NAND2_X1 U9285 ( .A1(n8012), .A2(n8011), .ZN(n8014) );
  INV_X1 U9286 ( .A(n8020), .ZN(n8013) );
  XNOR2_X1 U9287 ( .A(n8014), .B(n8013), .ZN(n8018) );
  OR2_X1 U9288 ( .A1(n8181), .A2(n10462), .ZN(n8017) );
  OR2_X1 U9289 ( .A1(n8015), .A2(n10464), .ZN(n8016) );
  NAND2_X1 U9290 ( .A1(n8017), .A2(n8016), .ZN(n8076) );
  AOI21_X1 U9291 ( .B1(n8018), .B2(n10821), .A(n8076), .ZN(n10842) );
  XNOR2_X1 U9292 ( .A(n8020), .B(n8019), .ZN(n10840) );
  NAND2_X1 U9293 ( .A1(n10814), .A2(n8072), .ZN(n8021) );
  NAND2_X1 U9294 ( .A1(n8021), .A2(n10949), .ZN(n8023) );
  OR2_X1 U9295 ( .A1(n8023), .A2(n8022), .ZN(n10837) );
  AOI22_X1 U9296 ( .A1(n11005), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n8079), .B2(
        n10992), .ZN(n8025) );
  NAND2_X1 U9297 ( .A1(n10956), .A2(n8072), .ZN(n8024) );
  OAI211_X1 U9298 ( .C1(n10837), .C2(n10477), .A(n8025), .B(n8024), .ZN(n8026)
         );
  AOI21_X1 U9299 ( .B1(n10840), .B2(n10961), .A(n8026), .ZN(n8027) );
  OAI21_X1 U9300 ( .B1(n10842), .B2(n11005), .A(n8027), .ZN(P1_U3288) );
  XNOR2_X1 U9301 ( .A(n8032), .B(n8028), .ZN(n8030) );
  OAI21_X1 U9302 ( .B1(n8030), .B2(n10941), .A(n8029), .ZN(n10805) );
  INV_X1 U9303 ( .A(n10805), .ZN(n8039) );
  XNOR2_X1 U9304 ( .A(n8031), .B(n8032), .ZN(n10807) );
  OAI211_X1 U9305 ( .C1(n10785), .C2(n7806), .A(n10813), .B(n10949), .ZN(
        n10803) );
  AOI22_X1 U9306 ( .A1(n11005), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10992), .B2(
        n8033), .ZN(n8036) );
  NAND2_X1 U9307 ( .A1(n10956), .A2(n8034), .ZN(n8035) );
  OAI211_X1 U9308 ( .C1(n10803), .C2(n10477), .A(n8036), .B(n8035), .ZN(n8037)
         );
  AOI21_X1 U9309 ( .B1(n10807), .B2(n10961), .A(n8037), .ZN(n8038) );
  OAI21_X1 U9310 ( .B1(n8039), .B2(n11005), .A(n8038), .ZN(P1_U3290) );
  INV_X1 U9311 ( .A(n8040), .ZN(n8043) );
  OAI222_X1 U9312 ( .A1(n8793), .A2(n8041), .B1(n8791), .B2(n8043), .C1(
        P1_U3086), .C2(n10219), .ZN(P1_U3336) );
  OAI222_X1 U9313 ( .A1(n9261), .A2(n8044), .B1(n9792), .B2(n8043), .C1(n8042), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  XNOR2_X1 U9314 ( .A(n8514), .B(n7766), .ZN(n8047) );
  NAND2_X1 U9315 ( .A1(n8047), .A2(n9397), .ZN(n8109) );
  NAND2_X1 U9316 ( .A1(n5185), .A2(n8109), .ZN(n8048) );
  XNOR2_X1 U9317 ( .A(n8110), .B(n8048), .ZN(n8054) );
  NOR2_X1 U9318 ( .A1(n9328), .A2(n8449), .ZN(n8049) );
  AOI211_X1 U9319 ( .C1(n9330), .C2(n9398), .A(n8050), .B(n8049), .ZN(n8051)
         );
  OAI21_X1 U9320 ( .B1(n5707), .B2(n9377), .A(n8051), .ZN(n8052) );
  AOI21_X1 U9321 ( .B1(n8452), .B2(n9353), .A(n8052), .ZN(n8053) );
  OAI21_X1 U9322 ( .B1(n8054), .B2(n9355), .A(n8053), .ZN(P2_U3161) );
  AOI21_X1 U9323 ( .B1(n8057), .B2(n8056), .A(n8055), .ZN(n8063) );
  NOR2_X1 U9324 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9116), .ZN(n10701) );
  OAI22_X1 U9325 ( .A1(n9376), .A2(n8058), .B1(n8349), .B2(n9383), .ZN(n8059)
         );
  AOI211_X1 U9326 ( .C1(n9380), .C2(n9399), .A(n10701), .B(n8059), .ZN(n8062)
         );
  INV_X1 U9327 ( .A(n8348), .ZN(n8060) );
  NAND2_X1 U9328 ( .A1(n9364), .A2(n8060), .ZN(n8061) );
  OAI211_X1 U9329 ( .C1(n8063), .C2(n9355), .A(n8062), .B(n8061), .ZN(P2_U3167) );
  OAI22_X1 U9330 ( .A1(n8071), .A2(n7808), .B1(n10838), .B2(n9860), .ZN(n8066)
         );
  XNOR2_X1 U9331 ( .A(n8066), .B(n9951), .ZN(n8069) );
  INV_X1 U9332 ( .A(n8069), .ZN(n8067) );
  NAND2_X1 U9333 ( .A1(n8147), .A2(n8146), .ZN(n8075) );
  OR2_X1 U9334 ( .A1(n8071), .A2(n9901), .ZN(n8074) );
  NAND2_X1 U9335 ( .A1(n8072), .A2(n9954), .ZN(n8073) );
  AND2_X1 U9336 ( .A1(n8074), .A2(n8073), .ZN(n8145) );
  XNOR2_X1 U9337 ( .A(n8075), .B(n8145), .ZN(n8081) );
  AOI22_X1 U9338 ( .A1(n8076), .A2(n10029), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3086), .ZN(n8077) );
  OAI21_X1 U9339 ( .B1(n10838), .B2(n10090), .A(n8077), .ZN(n8078) );
  AOI21_X1 U9340 ( .B1(n8079), .B2(n10071), .A(n8078), .ZN(n8080) );
  OAI21_X1 U9341 ( .B1(n8081), .B2(n10064), .A(n8080), .ZN(P1_U3227) );
  NAND2_X1 U9342 ( .A1(n8106), .A2(n10582), .ZN(n8083) );
  OAI211_X1 U9343 ( .C1(n8084), .C2(n8793), .A(n8083), .B(n8082), .ZN(P1_U3335) );
  INV_X1 U9344 ( .A(n8111), .ZN(n8480) );
  XNOR2_X1 U9345 ( .A(n8085), .B(n8086), .ZN(n8479) );
  OAI211_X1 U9346 ( .C1(n8088), .C2(n6205), .A(n9664), .B(n8087), .ZN(n8090)
         );
  AOI22_X1 U9347 ( .A1(n9396), .A2(n9668), .B1(n9667), .B2(n9397), .ZN(n8089)
         );
  NAND2_X1 U9348 ( .A1(n8090), .A2(n8089), .ZN(n8484) );
  AOI21_X1 U9349 ( .B1(n8479), .B2(n9733), .A(n8484), .ZN(n8092) );
  MUX2_X1 U9350 ( .A(n8138), .B(n8092), .S(n9735), .Z(n8091) );
  OAI21_X1 U9351 ( .B1(n8480), .B2(n9738), .A(n8091), .ZN(P2_U3468) );
  MUX2_X1 U9352 ( .A(n6198), .B(n8092), .S(n11017), .Z(n8093) );
  OAI21_X1 U9353 ( .B1(n8480), .B2(n9779), .A(n8093), .ZN(P2_U3417) );
  NAND2_X1 U9354 ( .A1(n8094), .A2(n8101), .ZN(n8095) );
  NAND2_X1 U9355 ( .A1(n8096), .A2(n8095), .ZN(n8099) );
  NAND2_X1 U9356 ( .A1(n9395), .A2(n9668), .ZN(n8097) );
  OAI21_X1 U9357 ( .B1(n8449), .B2(n9635), .A(n8097), .ZN(n8098) );
  AOI21_X1 U9358 ( .B1(n8099), .B2(n9664), .A(n8098), .ZN(n8296) );
  INV_X1 U9359 ( .A(n8101), .ZN(n8102) );
  XNOR2_X1 U9360 ( .A(n8100), .B(n8102), .ZN(n8293) );
  NAND2_X1 U9361 ( .A1(n8293), .A2(n9733), .ZN(n8104) );
  NAND2_X1 U9362 ( .A1(n8290), .A2(n9720), .ZN(n8103) );
  OR2_X1 U9363 ( .A1(n9735), .A2(n6214), .ZN(n8105) );
  OAI21_X1 U9364 ( .B1(n10923), .B2(n9683), .A(n8105), .ZN(P2_U3469) );
  INV_X1 U9365 ( .A(n8106), .ZN(n8107) );
  OAI222_X1 U9366 ( .A1(n9261), .A2(n8108), .B1(n9792), .B2(n8107), .C1(n6481), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  XNOR2_X1 U9367 ( .A(n8111), .B(n8831), .ZN(n8251) );
  XNOR2_X1 U9368 ( .A(n8251), .B(n8449), .ZN(n8112) );
  OAI211_X1 U9369 ( .C1(n8113), .C2(n8112), .A(n8254), .B(n5658), .ZN(n8119)
         );
  INV_X1 U9370 ( .A(n8481), .ZN(n8117) );
  NOR2_X1 U9371 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8114), .ZN(n8133) );
  AOI21_X1 U9372 ( .B1(n9330), .B2(n9397), .A(n8133), .ZN(n8115) );
  OAI21_X1 U9373 ( .B1(n8325), .B2(n9328), .A(n8115), .ZN(n8116) );
  AOI21_X1 U9374 ( .B1(n8117), .B2(n9364), .A(n8116), .ZN(n8118) );
  OAI211_X1 U9375 ( .C1(n8480), .C2(n9383), .A(n8119), .B(n8118), .ZN(P2_U3171) );
  INV_X1 U9376 ( .A(n8120), .ZN(n8124) );
  OAI222_X1 U9377 ( .A1(n9792), .A2(n8124), .B1(P2_U3151), .B2(n8122), .C1(
        n8121), .C2(n9783), .ZN(P2_U3274) );
  OAI222_X1 U9378 ( .A1(n8793), .A2(n8125), .B1(n8791), .B2(n8124), .C1(n8123), 
        .C2(P1_U3086), .ZN(P1_U3334) );
  AOI21_X1 U9379 ( .B1(n8128), .B2(n8127), .A(n8126), .ZN(n8144) );
  NAND2_X1 U9380 ( .A1(n8130), .A2(n8129), .ZN(n8131) );
  XNOR2_X1 U9381 ( .A(n8132), .B(n8131), .ZN(n8142) );
  AOI21_X1 U9382 ( .B1(n9505), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8133), .ZN(
        n8134) );
  OAI21_X1 U9383 ( .B1(n8135), .B2(n9521), .A(n8134), .ZN(n8141) );
  AOI21_X1 U9384 ( .B1(n8138), .B2(n8137), .A(n8136), .ZN(n8139) );
  NOR2_X1 U9385 ( .A1(n8139), .A2(n10717), .ZN(n8140) );
  AOI211_X1 U9386 ( .C1(n10729), .C2(n8142), .A(n8141), .B(n8140), .ZN(n8143)
         );
  OAI21_X1 U9387 ( .B1(n8144), .B2(n10724), .A(n8143), .ZN(P2_U3191) );
  OAI22_X1 U9388 ( .A1(n8181), .A2(n7808), .B1(n8002), .B2(n9860), .ZN(n8148)
         );
  XNOR2_X1 U9389 ( .A(n8148), .B(n9899), .ZN(n8153) );
  OR2_X1 U9390 ( .A1(n8181), .A2(n9901), .ZN(n8151) );
  NAND2_X1 U9391 ( .A1(n8149), .A2(n9954), .ZN(n8150) );
  NAND2_X1 U9392 ( .A1(n8151), .A2(n8150), .ZN(n8154) );
  INV_X1 U9393 ( .A(n8154), .ZN(n8152) );
  NAND2_X1 U9394 ( .A1(n8153), .A2(n8152), .ZN(n8161) );
  INV_X1 U9395 ( .A(n8153), .ZN(n8155) );
  NAND2_X1 U9396 ( .A1(n8155), .A2(n8154), .ZN(n8157) );
  INV_X1 U9397 ( .A(n8299), .ZN(n8162) );
  INV_X1 U9398 ( .A(n8156), .ZN(n8158) );
  NAND2_X1 U9399 ( .A1(n8158), .A2(n8157), .ZN(n8160) );
  AOI22_X1 U9400 ( .A1(n8162), .A2(n8161), .B1(n8160), .B2(n8159), .ZN(n8168)
         );
  AOI22_X1 U9401 ( .A1(n8163), .A2(n10029), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n8164) );
  OAI21_X1 U9402 ( .B1(n8002), .B2(n10090), .A(n8164), .ZN(n8165) );
  AOI21_X1 U9403 ( .B1(n8166), .B2(n10071), .A(n8165), .ZN(n8167) );
  OAI21_X1 U9404 ( .B1(n8168), .B2(n10064), .A(n8167), .ZN(P1_U3239) );
  NAND2_X1 U9405 ( .A1(n10099), .A2(n9953), .ZN(n8170) );
  OR2_X1 U9406 ( .A1(n10858), .A2(n7808), .ZN(n8169) );
  NAND2_X1 U9407 ( .A1(n8170), .A2(n8169), .ZN(n8298) );
  NAND2_X1 U9408 ( .A1(n10099), .A2(n9954), .ZN(n8172) );
  OR2_X1 U9409 ( .A1(n10858), .A2(n9860), .ZN(n8171) );
  NAND2_X1 U9410 ( .A1(n8172), .A2(n8171), .ZN(n8173) );
  XNOR2_X1 U9411 ( .A(n8173), .B(n9951), .ZN(n8297) );
  XOR2_X1 U9412 ( .A(n8298), .B(n8297), .Z(n8174) );
  XNOR2_X1 U9413 ( .A(n8299), .B(n8174), .ZN(n8178) );
  OAI22_X1 U9414 ( .A1(n8181), .A2(n10464), .B1(n8303), .B2(n10462), .ZN(n8187) );
  AOI22_X1 U9415 ( .A1(n8187), .A2(n10029), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n8175) );
  OAI21_X1 U9416 ( .B1(n8190), .B2(n10084), .A(n8175), .ZN(n8176) );
  AOI21_X1 U9417 ( .B1(n8192), .B2(n10073), .A(n8176), .ZN(n8177) );
  OAI21_X1 U9418 ( .B1(n8178), .B2(n10064), .A(n8177), .ZN(P1_U3213) );
  NAND2_X1 U9419 ( .A1(n8180), .A2(n8179), .ZN(n8183) );
  NAND2_X1 U9420 ( .A1(n8181), .A2(n8002), .ZN(n8182) );
  NAND2_X1 U9421 ( .A1(n8183), .A2(n8182), .ZN(n8273) );
  XNOR2_X1 U9422 ( .A(n8273), .B(n8186), .ZN(n10855) );
  INV_X1 U9423 ( .A(n8184), .ZN(n8185) );
  NOR2_X1 U9424 ( .A1(n8185), .A2(n8272), .ZN(n10887) );
  INV_X1 U9425 ( .A(n10887), .ZN(n10883) );
  OAI21_X1 U9426 ( .B1(n8184), .B2(n8186), .A(n10883), .ZN(n8188) );
  AOI21_X1 U9427 ( .B1(n8188), .B2(n10821), .A(n8187), .ZN(n10857) );
  INV_X1 U9428 ( .A(n10857), .ZN(n8196) );
  NAND2_X1 U9429 ( .A1(n8189), .A2(n10858), .ZN(n10878) );
  OAI211_X1 U9430 ( .C1(n8189), .C2(n10858), .A(n10949), .B(n10878), .ZN(
        n10856) );
  NOR2_X1 U9431 ( .A1(n10472), .A2(n8190), .ZN(n8191) );
  AOI21_X1 U9432 ( .B1(n11005), .B2(P1_REG2_REG_7__SCAN_IN), .A(n8191), .ZN(
        n8194) );
  NAND2_X1 U9433 ( .A1(n10956), .A2(n8192), .ZN(n8193) );
  OAI211_X1 U9434 ( .C1(n10856), .C2(n10477), .A(n8194), .B(n8193), .ZN(n8195)
         );
  AOI21_X1 U9435 ( .B1(n8196), .B2(n10475), .A(n8195), .ZN(n8197) );
  OAI21_X1 U9436 ( .B1(n10458), .B2(n10855), .A(n8197), .ZN(P1_U3286) );
  AOI21_X1 U9437 ( .B1(n8200), .B2(n8199), .A(n8198), .ZN(n8214) );
  INV_X1 U9438 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8206) );
  OAI21_X1 U9439 ( .B1(n8203), .B2(n8202), .A(n8201), .ZN(n8204) );
  NAND2_X1 U9440 ( .A1(n8204), .A2(n10729), .ZN(n8205) );
  NAND2_X1 U9441 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8255) );
  OAI211_X1 U9442 ( .C1(n10734), .C2(n8206), .A(n8205), .B(n8255), .ZN(n8211)
         );
  AOI21_X1 U9443 ( .B1(n8208), .B2(n8207), .A(n5181), .ZN(n8209) );
  NOR2_X1 U9444 ( .A1(n8209), .A2(n10724), .ZN(n8210) );
  AOI211_X1 U9445 ( .C1(n10722), .C2(n8212), .A(n8211), .B(n8210), .ZN(n8213)
         );
  OAI21_X1 U9446 ( .B1(n8214), .B2(n10717), .A(n8213), .ZN(P2_U3192) );
  INV_X1 U9447 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n8376) );
  MUX2_X1 U9448 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n8376), .S(n10105), .Z(
        n10112) );
  OAI21_X1 U9449 ( .B1(n8220), .B2(P1_REG2_REG_9__SCAN_IN), .A(n8215), .ZN(
        n8216) );
  NAND2_X1 U9450 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n8390), .ZN(n8217) );
  OAI21_X1 U9451 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n8390), .A(n8217), .ZN(
        n8218) );
  NOR2_X1 U9452 ( .A1(n8219), .A2(n8218), .ZN(n8389) );
  AOI211_X1 U9453 ( .C1(n8219), .C2(n8218), .A(n8389), .B(n10763), .ZN(n8232)
         );
  INV_X1 U9454 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10933) );
  MUX2_X1 U9455 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10933), .S(n8390), .Z(n8225) );
  INV_X1 U9456 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10920) );
  MUX2_X1 U9457 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n10920), .S(n10105), .Z(
        n10115) );
  OR2_X1 U9458 ( .A1(n8220), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8222) );
  NAND2_X1 U9459 ( .A1(n10115), .A2(n10114), .ZN(n10113) );
  NAND2_X1 U9460 ( .A1(n10105), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8223) );
  NAND2_X1 U9461 ( .A1(n10113), .A2(n8223), .ZN(n8224) );
  NAND2_X1 U9462 ( .A1(n8224), .A2(n8225), .ZN(n8384) );
  OAI211_X1 U9463 ( .C1(n8225), .C2(n8224), .A(n10147), .B(n8384), .ZN(n8226)
         );
  INV_X1 U9464 ( .A(n8226), .ZN(n8231) );
  INV_X1 U9465 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n8229) );
  NAND2_X1 U9466 ( .A1(n10770), .A2(n8390), .ZN(n8228) );
  NAND2_X1 U9467 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n8227) );
  OAI211_X1 U9468 ( .C1(n8229), .C2(n10203), .A(n8228), .B(n8227), .ZN(n8230)
         );
  OR3_X1 U9469 ( .A1(n8232), .A2(n8231), .A3(n8230), .ZN(P1_U3254) );
  INV_X1 U9470 ( .A(n8233), .ZN(n8234) );
  NAND2_X1 U9471 ( .A1(n8235), .A2(n8234), .ZN(n8240) );
  INV_X1 U9472 ( .A(n8236), .ZN(n8237) );
  NAND2_X1 U9473 ( .A1(n8238), .A2(n8237), .ZN(n8239) );
  NAND2_X1 U9474 ( .A1(n8240), .A2(n8239), .ZN(n8241) );
  NAND2_X1 U9475 ( .A1(n8242), .A2(n8241), .ZN(n8358) );
  AND2_X1 U9476 ( .A1(n8243), .A2(n7730), .ZN(n8291) );
  AND2_X1 U9477 ( .A1(n10874), .A2(n8291), .ZN(n9544) );
  OAI22_X1 U9478 ( .A1(n9647), .A2(n8245), .B1(n8244), .B2(n9590), .ZN(n8248)
         );
  MUX2_X1 U9479 ( .A(n8246), .B(P2_REG2_REG_1__SCAN_IN), .S(n9673), .Z(n8247)
         );
  AOI211_X1 U9480 ( .C1(n9544), .C2(n8249), .A(n8248), .B(n8247), .ZN(n8250)
         );
  INV_X1 U9481 ( .A(n8250), .ZN(P2_U3232) );
  NAND2_X1 U9482 ( .A1(n8251), .A2(n8252), .ZN(n8253) );
  NAND2_X1 U9483 ( .A1(n8254), .A2(n8253), .ZN(n8436) );
  XNOR2_X1 U9484 ( .A(n8290), .B(n7735), .ZN(n8435) );
  XNOR2_X1 U9485 ( .A(n8436), .B(n8435), .ZN(n8437) );
  XNOR2_X1 U9486 ( .A(n8437), .B(n8325), .ZN(n8260) );
  OAI21_X1 U9487 ( .B1(n9328), .B2(n8473), .A(n8255), .ZN(n8256) );
  AOI21_X1 U9488 ( .B1(n9330), .B2(n8252), .A(n8256), .ZN(n8257) );
  OAI21_X1 U9489 ( .B1(n9377), .B2(n8287), .A(n8257), .ZN(n8258) );
  AOI21_X1 U9490 ( .B1(n8290), .B2(n9353), .A(n8258), .ZN(n8259) );
  OAI21_X1 U9491 ( .B1(n8260), .B2(n9355), .A(n8259), .ZN(P2_U3157) );
  INV_X1 U9492 ( .A(n8261), .ZN(n8263) );
  OAI222_X1 U9493 ( .A1(n8793), .A2(n9156), .B1(n8791), .B2(n8263), .C1(
        P1_U3086), .C2(n5452), .ZN(P1_U3333) );
  OAI222_X1 U9494 ( .A1(n9261), .A2(n8264), .B1(n9792), .B2(n8263), .C1(n8262), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  XNOR2_X1 U9495 ( .A(n8265), .B(n8266), .ZN(n8267) );
  OAI222_X1 U9496 ( .A1(n9637), .A2(n8713), .B1(n9635), .B2(n8473), .C1(n8267), 
        .C2(n9653), .ZN(n8521) );
  XNOR2_X1 U9497 ( .A(n8268), .B(n6454), .ZN(n8527) );
  OAI22_X1 U9498 ( .A1(n8527), .A2(n9718), .B1(n8471), .B2(n8726), .ZN(n8269)
         );
  NOR2_X1 U9499 ( .A1(n8521), .A2(n8269), .ZN(n10936) );
  OR2_X1 U9500 ( .A1(n9735), .A2(n8270), .ZN(n8271) );
  OAI21_X1 U9501 ( .B1(n10936), .B2(n9683), .A(n8271), .ZN(P2_U3471) );
  NAND2_X1 U9502 ( .A1(n5344), .A2(n10858), .ZN(n8274) );
  NAND2_X1 U9503 ( .A1(n8275), .A2(n10884), .ZN(n10890) );
  NAND2_X1 U9504 ( .A1(n8277), .A2(n8276), .ZN(n8370) );
  XNOR2_X1 U9505 ( .A(n8371), .B(n8370), .ZN(n10911) );
  INV_X1 U9506 ( .A(n10911), .ZN(n8286) );
  OAI21_X1 U9507 ( .B1(n10887), .B2(n10885), .A(n10884), .ZN(n8278) );
  XOR2_X1 U9508 ( .A(n8370), .B(n8278), .Z(n8279) );
  OR2_X1 U9509 ( .A1(n8303), .A2(n10464), .ZN(n8339) );
  OAI21_X1 U9510 ( .B1(n8279), .B2(n10941), .A(n8339), .ZN(n10909) );
  AOI211_X1 U9511 ( .C1(n8345), .C2(n10879), .A(n10976), .B(n8378), .ZN(n8281)
         );
  NAND2_X1 U9512 ( .A1(n10096), .A2(n10552), .ZN(n8338) );
  INV_X1 U9513 ( .A(n8338), .ZN(n8280) );
  NOR2_X1 U9514 ( .A1(n8281), .A2(n8280), .ZN(n10907) );
  AOI22_X1 U9515 ( .A1(n11005), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8337), .B2(
        n10992), .ZN(n8283) );
  NAND2_X1 U9516 ( .A1(n10956), .A2(n8345), .ZN(n8282) );
  OAI211_X1 U9517 ( .C1(n10907), .C2(n10477), .A(n8283), .B(n8282), .ZN(n8284)
         );
  AOI21_X1 U9518 ( .B1(n10909), .B2(n10475), .A(n8284), .ZN(n8285) );
  OAI21_X1 U9519 ( .B1(n10458), .B2(n8286), .A(n8285), .ZN(P1_U3284) );
  INV_X2 U9520 ( .A(n9673), .ZN(n10874) );
  INV_X1 U9521 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8288) );
  OAI22_X1 U9522 ( .A1(n10874), .A2(n8288), .B1(n8287), .B2(n9590), .ZN(n8289)
         );
  AOI21_X1 U9523 ( .B1(n10869), .B2(n8290), .A(n8289), .ZN(n8295) );
  OR2_X1 U9524 ( .A1(n8292), .A2(n8291), .ZN(n10865) );
  NAND2_X1 U9525 ( .A1(n8293), .A2(n9677), .ZN(n8294) );
  OAI211_X1 U9526 ( .C1(n8296), .C2(n9673), .A(n8295), .B(n8294), .ZN(P2_U3223) );
  NAND2_X1 U9527 ( .A1(n8299), .A2(n8298), .ZN(n8300) );
  NAND2_X1 U9528 ( .A1(n8301), .A2(n8300), .ZN(n8329) );
  OAI22_X1 U9529 ( .A1(n8303), .A2(n7808), .B1(n10881), .B2(n9860), .ZN(n8302)
         );
  XNOR2_X1 U9530 ( .A(n8302), .B(n9899), .ZN(n8330) );
  OR2_X1 U9531 ( .A1(n8303), .A2(n9901), .ZN(n8305) );
  NAND2_X1 U9532 ( .A1(n10899), .A2(n9954), .ZN(n8304) );
  NAND2_X1 U9533 ( .A1(n8305), .A2(n8304), .ZN(n8331) );
  XNOR2_X1 U9534 ( .A(n8330), .B(n8331), .ZN(n8328) );
  XNOR2_X1 U9535 ( .A(n8329), .B(n8328), .ZN(n8310) );
  INV_X1 U9536 ( .A(n10898), .ZN(n8307) );
  OAI22_X1 U9537 ( .A1(n5344), .A2(n10464), .B1(n8372), .B2(n10462), .ZN(
        n10892) );
  AOI22_X1 U9538 ( .A1(n10892), .A2(n10029), .B1(P1_REG3_REG_8__SCAN_IN), .B2(
        P1_U3086), .ZN(n8306) );
  OAI21_X1 U9539 ( .B1(n8307), .B2(n10084), .A(n8306), .ZN(n8308) );
  AOI21_X1 U9540 ( .B1(n10899), .B2(n10073), .A(n8308), .ZN(n8309) );
  OAI21_X1 U9541 ( .B1(n8310), .B2(n10064), .A(n8309), .ZN(P1_U3221) );
  OAI22_X1 U9542 ( .A1(n9647), .A2(n8312), .B1(n8311), .B2(n9590), .ZN(n8315)
         );
  MUX2_X1 U9543 ( .A(n8313), .B(P2_REG2_REG_4__SCAN_IN), .S(n9673), .Z(n8314)
         );
  AOI211_X1 U9544 ( .C1(n9677), .C2(n8316), .A(n8315), .B(n8314), .ZN(n8317)
         );
  INV_X1 U9545 ( .A(n8317), .ZN(P2_U3229) );
  INV_X1 U9546 ( .A(n8318), .ZN(n8319) );
  AOI21_X1 U9547 ( .B1(n8100), .B2(n8320), .A(n8319), .ZN(n8321) );
  XOR2_X1 U9548 ( .A(n8322), .B(n8321), .Z(n8547) );
  NOR2_X1 U9549 ( .A1(n8547), .A2(n9718), .ZN(n8326) );
  XNOR2_X1 U9550 ( .A(n8323), .B(n8322), .ZN(n8324) );
  OAI222_X1 U9551 ( .A1(n9635), .A2(n8325), .B1(n9637), .B2(n8660), .C1(n8324), 
        .C2(n9653), .ZN(n8541) );
  AOI211_X1 U9552 ( .C1(n9720), .C2(n8544), .A(n8326), .B(n8541), .ZN(n10924)
         );
  NAND2_X1 U9553 ( .A1(n9683), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8327) );
  OAI21_X1 U9554 ( .B1(n10924), .B2(n9683), .A(n8327), .ZN(P2_U3470) );
  INV_X1 U9555 ( .A(n8330), .ZN(n8332) );
  NAND2_X1 U9556 ( .A1(n8332), .A2(n8331), .ZN(n8333) );
  OAI22_X1 U9557 ( .A1(n8372), .A2(n7808), .B1(n10908), .B2(n9860), .ZN(n8334)
         );
  XNOR2_X1 U9558 ( .A(n8334), .B(n9899), .ZN(n8567) );
  OR2_X1 U9559 ( .A1(n8372), .A2(n9901), .ZN(n8336) );
  NAND2_X1 U9560 ( .A1(n8345), .A2(n9954), .ZN(n8335) );
  NAND2_X1 U9561 ( .A1(n8336), .A2(n8335), .ZN(n8568) );
  XNOR2_X1 U9562 ( .A(n8567), .B(n8568), .ZN(n8565) );
  XNOR2_X1 U9563 ( .A(n8566), .B(n8565), .ZN(n8347) );
  INV_X1 U9564 ( .A(n8337), .ZN(n8343) );
  NAND2_X1 U9565 ( .A1(n8339), .A2(n8338), .ZN(n8340) );
  NAND2_X1 U9566 ( .A1(n8340), .A2(n10029), .ZN(n8342) );
  OAI211_X1 U9567 ( .C1(n10084), .C2(n8343), .A(n8342), .B(n8341), .ZN(n8344)
         );
  AOI21_X1 U9568 ( .B1(n8345), .B2(n10073), .A(n8344), .ZN(n8346) );
  OAI21_X1 U9569 ( .B1(n8347), .B2(n10064), .A(n8346), .ZN(P1_U3231) );
  OAI22_X1 U9570 ( .A1(n9647), .A2(n8349), .B1(n8348), .B2(n9590), .ZN(n8352)
         );
  MUX2_X1 U9571 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n8350), .S(n10874), .Z(n8351)
         );
  AOI211_X1 U9572 ( .C1(n9677), .C2(n8353), .A(n8352), .B(n8351), .ZN(n8354)
         );
  INV_X1 U9573 ( .A(n8354), .ZN(P2_U3228) );
  NAND3_X1 U9574 ( .A1(n8356), .A2(n8355), .A3(n8726), .ZN(n8359) );
  OAI22_X1 U9575 ( .A1(n8359), .A2(n8358), .B1(n8357), .B2(n9590), .ZN(n8362)
         );
  MUX2_X1 U9576 ( .A(P2_REG2_REG_0__SCAN_IN), .B(n8360), .S(n10874), .Z(n8361)
         );
  AOI211_X1 U9577 ( .C1(n10869), .C2(n8363), .A(n8362), .B(n8361), .ZN(n8364)
         );
  INV_X1 U9578 ( .A(n8364), .ZN(P2_U3233) );
  XNOR2_X1 U9579 ( .A(n8365), .B(n8366), .ZN(n8369) );
  OR2_X1 U9580 ( .A1(n8746), .A2(n10462), .ZN(n8368) );
  OR2_X1 U9581 ( .A1(n8372), .A2(n10464), .ZN(n8367) );
  NAND2_X1 U9582 ( .A1(n8368), .A2(n8367), .ZN(n8579) );
  AOI21_X1 U9583 ( .B1(n8369), .B2(n10821), .A(n8579), .ZN(n10916) );
  NAND2_X1 U9584 ( .A1(n8371), .A2(n8370), .ZN(n8374) );
  NAND2_X1 U9585 ( .A1(n8372), .A2(n10908), .ZN(n8373) );
  NAND2_X1 U9586 ( .A1(n8374), .A2(n8373), .ZN(n8426) );
  XNOR2_X1 U9587 ( .A(n8426), .B(n8425), .ZN(n10919) );
  NAND2_X1 U9588 ( .A1(n10919), .A2(n10961), .ZN(n8382) );
  INV_X1 U9589 ( .A(n8375), .ZN(n8581) );
  OAI22_X1 U9590 ( .A1(n10475), .A2(n8376), .B1(n8581), .B2(n10472), .ZN(n8380) );
  INV_X1 U9591 ( .A(n8430), .ZN(n8377) );
  OAI211_X1 U9592 ( .C1(n10917), .C2(n8378), .A(n8377), .B(n10949), .ZN(n10915) );
  NOR2_X1 U9593 ( .A1(n10915), .A2(n10477), .ZN(n8379) );
  AOI211_X1 U9594 ( .C1(n10956), .C2(n8583), .A(n8380), .B(n8379), .ZN(n8381)
         );
  OAI211_X1 U9595 ( .C1(n11005), .C2(n10916), .A(n8382), .B(n8381), .ZN(
        P1_U3283) );
  INV_X1 U9596 ( .A(n8594), .ZN(n8398) );
  NAND2_X1 U9597 ( .A1(n8390), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8383) );
  INV_X1 U9598 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n8385) );
  MUX2_X1 U9599 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n8385), .S(n8594), .Z(n8386)
         );
  NAND2_X1 U9600 ( .A1(n8386), .A2(n8387), .ZN(n8593) );
  OAI21_X1 U9601 ( .B1(n8387), .B2(n8386), .A(n8593), .ZN(n8394) );
  NOR2_X1 U9602 ( .A1(n8594), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n8388) );
  AOI21_X1 U9603 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n8594), .A(n8388), .ZN(
        n8392) );
  AOI21_X1 U9604 ( .B1(n8390), .B2(P1_REG2_REG_11__SCAN_IN), .A(n8389), .ZN(
        n8391) );
  NAND2_X1 U9605 ( .A1(n8392), .A2(n8391), .ZN(n8588) );
  OAI21_X1 U9606 ( .B1(n8392), .B2(n8391), .A(n8588), .ZN(n8393) );
  AOI22_X1 U9607 ( .A1(n10147), .A2(n8394), .B1(n10222), .B2(n8393), .ZN(n8397) );
  NAND2_X1 U9608 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n8749) );
  INV_X1 U9609 ( .A(n8749), .ZN(n8395) );
  AOI21_X1 U9610 ( .B1(n10756), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n8395), .ZN(
        n8396) );
  OAI211_X1 U9611 ( .C1(n8398), .C2(n10220), .A(n8397), .B(n8396), .ZN(
        P1_U3255) );
  INV_X1 U9612 ( .A(n8399), .ZN(n8406) );
  NOR2_X1 U9613 ( .A1(n10874), .A2(n8400), .ZN(n8403) );
  OAI22_X1 U9614 ( .A1(n9647), .A2(n8401), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9590), .ZN(n8402) );
  AOI211_X1 U9615 ( .C1(n8404), .C2(n9677), .A(n8403), .B(n8402), .ZN(n8405)
         );
  OAI21_X1 U9616 ( .B1(n8406), .B2(n9673), .A(n8405), .ZN(P2_U3230) );
  INV_X1 U9617 ( .A(n8407), .ZN(n8414) );
  NOR2_X1 U9618 ( .A1(n9647), .A2(n8408), .ZN(n8411) );
  OAI22_X1 U9619 ( .A1(n10874), .A2(n5826), .B1(n8409), .B2(n9590), .ZN(n8410)
         );
  AOI211_X1 U9620 ( .C1(n8412), .C2(n9677), .A(n8411), .B(n8410), .ZN(n8413)
         );
  OAI21_X1 U9621 ( .B1(n8414), .B2(n9673), .A(n8413), .ZN(P2_U3227) );
  NAND2_X1 U9622 ( .A1(n8418), .A2(n9787), .ZN(n8416) );
  OAI211_X1 U9623 ( .C1(n8417), .C2(n9261), .A(n8416), .B(n8415), .ZN(P2_U3272) );
  NAND2_X1 U9624 ( .A1(n8418), .A2(n10582), .ZN(n8420) );
  OAI211_X1 U9625 ( .C1(n9155), .C2(n8793), .A(n8420), .B(n8419), .ZN(P1_U3332) );
  AOI21_X1 U9626 ( .B1(n8421), .B2(n8555), .A(n10941), .ZN(n8424) );
  OR2_X1 U9627 ( .A1(n10094), .A2(n10462), .ZN(n8423) );
  NAND2_X1 U9628 ( .A1(n10096), .A2(n10550), .ZN(n8422) );
  NAND2_X1 U9629 ( .A1(n8423), .A2(n8422), .ZN(n8615) );
  AOI21_X1 U9630 ( .B1(n8424), .B2(n10943), .A(n8615), .ZN(n10926) );
  NAND2_X1 U9631 ( .A1(n10917), .A2(n8427), .ZN(n8428) );
  XOR2_X1 U9632 ( .A(n8556), .B(n8555), .Z(n10929) );
  INV_X1 U9633 ( .A(n10929), .ZN(n10932) );
  NAND2_X1 U9634 ( .A1(n10932), .A2(n10961), .ZN(n8434) );
  INV_X1 U9635 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n8429) );
  OAI22_X1 U9636 ( .A1(n10475), .A2(n8429), .B1(n8617), .B2(n10472), .ZN(n8432) );
  INV_X1 U9637 ( .A(n8619), .ZN(n10927) );
  OAI211_X1 U9638 ( .C1(n8430), .C2(n10927), .A(n10949), .B(n10947), .ZN(
        n10925) );
  NOR2_X1 U9639 ( .A1(n10925), .A2(n10477), .ZN(n8431) );
  AOI211_X1 U9640 ( .C1(n10956), .C2(n8619), .A(n8432), .B(n8431), .ZN(n8433)
         );
  OAI211_X1 U9641 ( .C1(n10955), .C2(n10926), .A(n8434), .B(n8433), .ZN(
        P1_U3282) );
  XNOR2_X1 U9642 ( .A(n8544), .B(n8831), .ZN(n8467) );
  XNOR2_X1 U9643 ( .A(n8467), .B(n8473), .ZN(n8469) );
  XOR2_X1 U9644 ( .A(n8469), .B(n8470), .Z(n8442) );
  NAND2_X1 U9645 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8501) );
  OAI21_X1 U9646 ( .B1(n9328), .B2(n8660), .A(n8501), .ZN(n8438) );
  AOI21_X1 U9647 ( .B1(n9330), .B2(n9396), .A(n8438), .ZN(n8439) );
  OAI21_X1 U9648 ( .B1(n9377), .B2(n8542), .A(n8439), .ZN(n8440) );
  AOI21_X1 U9649 ( .B1(n8544), .B2(n9353), .A(n8440), .ZN(n8441) );
  OAI21_X1 U9650 ( .B1(n8442), .B2(n9355), .A(n8441), .ZN(P2_U3176) );
  NAND2_X1 U9651 ( .A1(n7882), .A2(n8443), .ZN(n8444) );
  XNOR2_X1 U9652 ( .A(n8444), .B(n8447), .ZN(n8513) );
  XOR2_X1 U9653 ( .A(n8447), .B(n5179), .Z(n8448) );
  OAI222_X1 U9654 ( .A1(n9637), .A2(n8449), .B1(n9635), .B2(n5647), .C1(n9653), 
        .C2(n8448), .ZN(n8518) );
  AOI21_X1 U9655 ( .B1(n9733), .B2(n8513), .A(n8518), .ZN(n8455) );
  OAI22_X1 U9656 ( .A1(n9779), .A2(n8514), .B1(n11017), .B2(n6181), .ZN(n8450)
         );
  INV_X1 U9657 ( .A(n8450), .ZN(n8451) );
  OAI21_X1 U9658 ( .B1(n8455), .B2(n11015), .A(n8451), .ZN(P2_U3414) );
  AOI22_X1 U9659 ( .A1(n8453), .A2(n8452), .B1(n9683), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n8454) );
  OAI21_X1 U9660 ( .B1(n8455), .B2(n9683), .A(n8454), .ZN(P2_U3467) );
  INV_X1 U9661 ( .A(n8456), .ZN(n8457) );
  AOI21_X1 U9662 ( .B1(n8461), .B2(n8458), .A(n8457), .ZN(n8459) );
  OAI222_X1 U9663 ( .A1(n9637), .A2(n8767), .B1(n9635), .B2(n8660), .C1(n9653), 
        .C2(n8459), .ZN(n8654) );
  INV_X1 U9664 ( .A(n8654), .ZN(n8466) );
  OAI21_X1 U9665 ( .B1(n8462), .B2(n8461), .A(n8460), .ZN(n8656) );
  INV_X1 U9666 ( .A(n8658), .ZN(n8675) );
  NOR2_X1 U9667 ( .A1(n8675), .A2(n9647), .ZN(n8464) );
  OAI22_X1 U9668 ( .A1(n10874), .A2(n5568), .B1(n8668), .B2(n9590), .ZN(n8463)
         );
  AOI211_X1 U9669 ( .C1(n8656), .C2(n9677), .A(n8464), .B(n8463), .ZN(n8465)
         );
  OAI21_X1 U9670 ( .B1(n8466), .B2(n9673), .A(n8465), .ZN(P2_U3220) );
  INV_X1 U9671 ( .A(n8467), .ZN(n8468) );
  XNOR2_X1 U9672 ( .A(n8471), .B(n8831), .ZN(n8661) );
  XNOR2_X1 U9673 ( .A(n8661), .B(n9394), .ZN(n8472) );
  XNOR2_X1 U9674 ( .A(n8664), .B(n8472), .ZN(n8478) );
  NAND2_X1 U9675 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9413) );
  OAI21_X1 U9676 ( .B1(n9376), .B2(n8473), .A(n9413), .ZN(n8474) );
  AOI21_X1 U9677 ( .B1(n9380), .B2(n9393), .A(n8474), .ZN(n8475) );
  OAI21_X1 U9678 ( .B1(n8522), .B2(n9377), .A(n8475), .ZN(n8476) );
  AOI21_X1 U9679 ( .B1(n8524), .B2(n9353), .A(n8476), .ZN(n8477) );
  OAI21_X1 U9680 ( .B1(n8478), .B2(n9355), .A(n8477), .ZN(P2_U3164) );
  INV_X1 U9681 ( .A(n8479), .ZN(n8486) );
  NOR2_X1 U9682 ( .A1(n8480), .A2(n9647), .ZN(n8483) );
  OAI22_X1 U9683 ( .A1(n10874), .A2(n8127), .B1(n8481), .B2(n9590), .ZN(n8482)
         );
  AOI211_X1 U9684 ( .C1(n8484), .C2(n10874), .A(n8483), .B(n8482), .ZN(n8485)
         );
  OAI21_X1 U9685 ( .B1(n9629), .B2(n8486), .A(n8485), .ZN(P2_U3224) );
  INV_X1 U9686 ( .A(n8487), .ZN(n8494) );
  NOR2_X1 U9687 ( .A1(n9590), .A2(n8488), .ZN(n8490) );
  AOI211_X1 U9688 ( .C1(n8491), .C2(n7729), .A(n8490), .B(n8489), .ZN(n8492)
         );
  MUX2_X1 U9689 ( .A(n5818), .B(n8492), .S(n10874), .Z(n8493) );
  OAI21_X1 U9690 ( .B1(n9629), .B2(n8494), .A(n8493), .ZN(P2_U3231) );
  AOI21_X1 U9691 ( .B1(n8497), .B2(n8496), .A(n8495), .ZN(n8512) );
  AOI21_X1 U9692 ( .B1(n8500), .B2(n8499), .A(n8498), .ZN(n8503) );
  NAND2_X1 U9693 ( .A1(n9505), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n8502) );
  OAI211_X1 U9694 ( .C1(n8503), .C2(n10724), .A(n8502), .B(n8501), .ZN(n8504)
         );
  AOI21_X1 U9695 ( .B1(n8505), .B2(n10722), .A(n8504), .ZN(n8511) );
  OAI21_X1 U9696 ( .B1(n8508), .B2(n8507), .A(n8506), .ZN(n8509) );
  NAND2_X1 U9697 ( .A1(n8509), .A2(n10729), .ZN(n8510) );
  OAI211_X1 U9698 ( .C1(n8512), .C2(n10717), .A(n8511), .B(n8510), .ZN(
        P2_U3193) );
  INV_X1 U9699 ( .A(n8513), .ZN(n8520) );
  NOR2_X1 U9700 ( .A1(n9647), .A2(n8514), .ZN(n8517) );
  OAI22_X1 U9701 ( .A1(n10874), .A2(n8515), .B1(n5707), .B2(n9590), .ZN(n8516)
         );
  AOI211_X1 U9702 ( .C1(n8518), .C2(n10874), .A(n8517), .B(n8516), .ZN(n8519)
         );
  OAI21_X1 U9703 ( .B1(n8520), .B2(n9629), .A(n8519), .ZN(P2_U3225) );
  NAND2_X1 U9704 ( .A1(n8521), .A2(n10874), .ZN(n8526) );
  OAI22_X1 U9705 ( .A1(n10874), .A2(n5842), .B1(n8522), .B2(n9590), .ZN(n8523)
         );
  AOI21_X1 U9706 ( .B1(n8524), .B2(n10869), .A(n8523), .ZN(n8525) );
  OAI211_X1 U9707 ( .C1(n8527), .C2(n9629), .A(n8526), .B(n8525), .ZN(P2_U3221) );
  NOR2_X1 U9708 ( .A1(n8529), .A2(n5366), .ZN(n8531) );
  INV_X1 U9709 ( .A(n8530), .ZN(n8623) );
  AOI21_X1 U9710 ( .B1(n8531), .B2(n8460), .A(n8623), .ZN(n8690) );
  AND2_X1 U9711 ( .A1(n8456), .A2(n8532), .ZN(n8535) );
  OAI211_X1 U9712 ( .C1(n8535), .C2(n8534), .A(n8533), .B(n9664), .ZN(n8537)
         );
  OR2_X1 U9713 ( .A1(n8713), .A2(n9635), .ZN(n8536) );
  OAI211_X1 U9714 ( .C1(n9307), .C2(n9637), .A(n8537), .B(n8536), .ZN(n8691)
         );
  NAND2_X1 U9715 ( .A1(n8691), .A2(n10874), .ZN(n8540) );
  OAI22_X1 U9716 ( .A1(n10874), .A2(n5847), .B1(n8714), .B2(n9590), .ZN(n8538)
         );
  AOI21_X1 U9717 ( .B1(n8706), .B2(n10869), .A(n8538), .ZN(n8539) );
  OAI211_X1 U9718 ( .C1(n8690), .C2(n9629), .A(n8540), .B(n8539), .ZN(P2_U3219) );
  NAND2_X1 U9719 ( .A1(n8541), .A2(n10874), .ZN(n8546) );
  OAI22_X1 U9720 ( .A1(n10874), .A2(n8499), .B1(n8542), .B2(n9590), .ZN(n8543)
         );
  AOI21_X1 U9721 ( .B1(n8544), .B2(n10869), .A(n8543), .ZN(n8545) );
  OAI211_X1 U9722 ( .C1(n8547), .C2(n9629), .A(n8546), .B(n8545), .ZN(P2_U3222) );
  NAND2_X1 U9723 ( .A1(n10946), .A2(n8548), .ZN(n8549) );
  NAND2_X1 U9724 ( .A1(n8549), .A2(n8635), .ZN(n8551) );
  NAND2_X1 U9725 ( .A1(n8551), .A2(n8550), .ZN(n8554) );
  OR2_X1 U9726 ( .A1(n10094), .A2(n10464), .ZN(n8553) );
  NAND2_X1 U9727 ( .A1(n10551), .A2(n10552), .ZN(n8552) );
  NAND2_X1 U9728 ( .A1(n8553), .A2(n8552), .ZN(n10039) );
  AOI21_X1 U9729 ( .B1(n8554), .B2(n10821), .A(n10039), .ZN(n10967) );
  NAND2_X1 U9730 ( .A1(n10937), .A2(n10938), .ZN(n8558) );
  INV_X1 U9731 ( .A(n10957), .ZN(n10950) );
  NAND2_X1 U9732 ( .A1(n10950), .A2(n10094), .ZN(n8557) );
  XNOR2_X1 U9733 ( .A(n8636), .B(n8635), .ZN(n10970) );
  NAND2_X1 U9734 ( .A1(n10970), .A2(n10961), .ZN(n8564) );
  INV_X1 U9735 ( .A(n9799), .ZN(n10968) );
  INV_X1 U9736 ( .A(n8644), .ZN(n8559) );
  OAI211_X1 U9737 ( .C1(n10968), .C2(n5405), .A(n8559), .B(n10949), .ZN(n10966) );
  INV_X1 U9738 ( .A(n10966), .ZN(n8562) );
  AOI22_X1 U9739 ( .A1(n11005), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n10044), 
        .B2(n10992), .ZN(n8560) );
  OAI21_X1 U9740 ( .B1(n10968), .B2(n10995), .A(n8560), .ZN(n8561) );
  AOI21_X1 U9741 ( .B1(n8562), .B2(n10959), .A(n8561), .ZN(n8563) );
  OAI211_X1 U9742 ( .C1(n11005), .C2(n10967), .A(n8564), .B(n8563), .ZN(
        P1_U3280) );
  INV_X1 U9743 ( .A(n8567), .ZN(n8569) );
  NAND2_X1 U9744 ( .A1(n10096), .A2(n9954), .ZN(n8570) );
  OAI21_X1 U9745 ( .B1(n10917), .B2(n9860), .A(n8570), .ZN(n8571) );
  XNOR2_X1 U9746 ( .A(n8571), .B(n9951), .ZN(n8574) );
  INV_X1 U9747 ( .A(n8574), .ZN(n8572) );
  NAND2_X1 U9748 ( .A1(n8604), .A2(n8603), .ZN(n8578) );
  OR2_X1 U9749 ( .A1(n10917), .A2(n7808), .ZN(n8577) );
  NAND2_X1 U9750 ( .A1(n10096), .A2(n9953), .ZN(n8576) );
  AND2_X1 U9751 ( .A1(n8577), .A2(n8576), .ZN(n8602) );
  XNOR2_X1 U9752 ( .A(n8578), .B(n8602), .ZN(n8585) );
  AOI22_X1 U9753 ( .A1(n8579), .A2(n10029), .B1(P1_REG3_REG_10__SCAN_IN), .B2(
        P1_U3086), .ZN(n8580) );
  OAI21_X1 U9754 ( .B1(n8581), .B2(n10084), .A(n8580), .ZN(n8582) );
  AOI21_X1 U9755 ( .B1(n8583), .B2(n10073), .A(n8582), .ZN(n8584) );
  OAI21_X1 U9756 ( .B1(n8585), .B2(n10064), .A(n8584), .ZN(P1_U3217) );
  INV_X1 U9757 ( .A(n8586), .ZN(n8677) );
  OAI222_X1 U9758 ( .A1(P1_U3086), .A2(n8587), .B1(n8791), .B2(n8677), .C1(
        n9154), .C2(n8793), .ZN(P1_U3331) );
  OAI21_X1 U9759 ( .B1(n8594), .B2(P1_REG2_REG_12__SCAN_IN), .A(n8588), .ZN(
        n8591) );
  NAND2_X1 U9760 ( .A1(n10124), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8589) );
  OAI21_X1 U9761 ( .B1(n10124), .B2(P1_REG2_REG_13__SCAN_IN), .A(n8589), .ZN(
        n8590) );
  AOI211_X1 U9762 ( .C1(n8591), .C2(n8590), .A(n10123), .B(n10763), .ZN(n8601)
         );
  INV_X1 U9763 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10971) );
  NOR2_X1 U9764 ( .A1(n10124), .A2(n10971), .ZN(n8592) );
  AOI21_X1 U9765 ( .B1(n10124), .B2(n10971), .A(n8592), .ZN(n8596) );
  OAI21_X1 U9766 ( .B1(n8594), .B2(P1_REG1_REG_12__SCAN_IN), .A(n8593), .ZN(
        n8595) );
  NOR2_X1 U9767 ( .A1(n8596), .A2(n8595), .ZN(n10127) );
  AOI211_X1 U9768 ( .C1(n8596), .C2(n8595), .A(n10127), .B(n10759), .ZN(n8600)
         );
  INV_X1 U9769 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U9770 ( .A1(n10770), .A2(n10124), .ZN(n8597) );
  NAND2_X1 U9771 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n10040) );
  OAI211_X1 U9772 ( .C1(n8598), .C2(n10203), .A(n8597), .B(n10040), .ZN(n8599)
         );
  OR3_X1 U9773 ( .A1(n8601), .A2(n8600), .A3(n8599), .ZN(P1_U3256) );
  NAND2_X1 U9774 ( .A1(n8603), .A2(n8602), .ZN(n8605) );
  NAND2_X1 U9775 ( .A1(n8619), .A2(n9948), .ZN(n8607) );
  OR2_X1 U9776 ( .A1(n8746), .A2(n7808), .ZN(n8606) );
  NAND2_X1 U9777 ( .A1(n8607), .A2(n8606), .ZN(n8608) );
  XNOR2_X1 U9778 ( .A(n8608), .B(n9899), .ZN(n8610) );
  AOI22_X1 U9779 ( .A1(n8619), .A2(n9954), .B1(n8609), .B2(n9953), .ZN(n8611)
         );
  INV_X1 U9780 ( .A(n8610), .ZN(n8613) );
  INV_X1 U9781 ( .A(n8611), .ZN(n8612) );
  NAND2_X1 U9782 ( .A1(n8613), .A2(n8612), .ZN(n8740) );
  NAND2_X1 U9783 ( .A1(n5711), .A2(n8740), .ZN(n8614) );
  XNOR2_X1 U9784 ( .A(n8739), .B(n8614), .ZN(n8621) );
  AOI22_X1 U9785 ( .A1(n8615), .A2(n10029), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n8616) );
  OAI21_X1 U9786 ( .B1(n8617), .B2(n10084), .A(n8616), .ZN(n8618) );
  AOI21_X1 U9787 ( .B1(n8619), .B2(n10073), .A(n8618), .ZN(n8620) );
  OAI21_X1 U9788 ( .B1(n8621), .B2(n10064), .A(n8620), .ZN(P1_U3236) );
  OAI21_X1 U9789 ( .B1(n8623), .B2(n8622), .A(n8626), .ZN(n8625) );
  NAND2_X1 U9790 ( .A1(n8625), .A2(n8624), .ZN(n8686) );
  XNOR2_X1 U9791 ( .A(n8627), .B(n8626), .ZN(n8628) );
  OAI222_X1 U9792 ( .A1(n9637), .A2(n8806), .B1(n9635), .B2(n8767), .C1(n8628), 
        .C2(n9653), .ZN(n8687) );
  NAND2_X1 U9793 ( .A1(n8687), .A2(n10874), .ZN(n8631) );
  OAI22_X1 U9794 ( .A1(n10874), .A2(n9468), .B1(n8768), .B2(n9590), .ZN(n8629)
         );
  AOI21_X1 U9795 ( .B1(n8760), .B2(n10869), .A(n8629), .ZN(n8630) );
  OAI211_X1 U9796 ( .C1(n8686), .C2(n9629), .A(n8631), .B(n8630), .ZN(P2_U3218) );
  INV_X1 U9797 ( .A(n8632), .ZN(n8652) );
  OAI222_X1 U9798 ( .A1(n9792), .A2(n8652), .B1(P2_U3151), .B2(n6485), .C1(
        n8633), .C2(n9783), .ZN(P2_U3270) );
  INV_X1 U9799 ( .A(n9924), .ZN(n10093) );
  NOR2_X1 U9800 ( .A1(n9799), .A2(n10093), .ZN(n8634) );
  INV_X1 U9801 ( .A(n8638), .ZN(n8637) );
  XNOR2_X1 U9802 ( .A(n10254), .B(n8637), .ZN(n10980) );
  XNOR2_X1 U9803 ( .A(n8639), .B(n8638), .ZN(n8642) );
  OAI22_X1 U9804 ( .A1(n9924), .A2(n10464), .B1(n10465), .B2(n10462), .ZN(
        n8640) );
  INV_X1 U9805 ( .A(n8640), .ZN(n8641) );
  OAI21_X1 U9806 ( .B1(n8642), .B2(n10941), .A(n8641), .ZN(n8643) );
  AOI21_X1 U9807 ( .B1(n10980), .B2(n10990), .A(n8643), .ZN(n10982) );
  INV_X1 U9808 ( .A(n10997), .ZN(n10902) );
  OR2_X1 U9809 ( .A1(n8644), .A2(n10975), .ZN(n8645) );
  NAND2_X1 U9810 ( .A1(n10555), .A2(n8645), .ZN(n10977) );
  INV_X1 U9811 ( .A(n11001), .ZN(n8648) );
  AOI22_X1 U9812 ( .A1(n11005), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9922), .B2(
        n10992), .ZN(n8647) );
  NAND2_X1 U9813 ( .A1(n10255), .A2(n10956), .ZN(n8646) );
  OAI211_X1 U9814 ( .C1(n10977), .C2(n8648), .A(n8647), .B(n8646), .ZN(n8649)
         );
  AOI21_X1 U9815 ( .B1(n10980), .B2(n10902), .A(n8649), .ZN(n8650) );
  OAI21_X1 U9816 ( .B1(n10982), .B2(n11005), .A(n8650), .ZN(P1_U3279) );
  OAI222_X1 U9817 ( .A1(P1_U3086), .A2(n8653), .B1(n8791), .B2(n8652), .C1(
        n8651), .C2(n8793), .ZN(P1_U3330) );
  NOR2_X1 U9818 ( .A1(n8675), .A2(n8726), .ZN(n8655) );
  AOI211_X1 U9819 ( .C1(n9733), .C2(n8656), .A(n8655), .B(n8654), .ZN(n10974)
         );
  OR2_X1 U9820 ( .A1(n10974), .A2(n9683), .ZN(n8657) );
  OAI21_X1 U9821 ( .B1(n9735), .B2(n9437), .A(n8657), .ZN(P2_U3472) );
  XNOR2_X1 U9822 ( .A(n8658), .B(n8831), .ZN(n8659) );
  NOR2_X1 U9823 ( .A1(n8659), .A2(n9393), .ZN(n8707) );
  AOI21_X1 U9824 ( .B1(n9393), .B2(n8659), .A(n8707), .ZN(n8666) );
  NAND2_X1 U9825 ( .A1(n8661), .A2(n8660), .ZN(n8663) );
  INV_X1 U9826 ( .A(n8661), .ZN(n8662) );
  OAI21_X1 U9827 ( .B1(n8666), .B2(n8665), .A(n8708), .ZN(n8667) );
  NAND2_X1 U9828 ( .A1(n8667), .A2(n5658), .ZN(n8674) );
  INV_X1 U9829 ( .A(n8668), .ZN(n8672) );
  NOR2_X1 U9830 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8669), .ZN(n9427) );
  AOI21_X1 U9831 ( .B1(n9330), .B2(n9394), .A(n9427), .ZN(n8670) );
  OAI21_X1 U9832 ( .B1(n8767), .B2(n9328), .A(n8670), .ZN(n8671) );
  AOI21_X1 U9833 ( .B1(n8672), .B2(n9364), .A(n8671), .ZN(n8673) );
  OAI211_X1 U9834 ( .C1(n8675), .C2(n9383), .A(n8674), .B(n8673), .ZN(P2_U3174) );
  OAI222_X1 U9835 ( .A1(n9792), .A2(n8677), .B1(P2_U3151), .B2(n6484), .C1(
        n8676), .C2(n9783), .ZN(P2_U3271) );
  XNOR2_X1 U9836 ( .A(n8679), .B(n8678), .ZN(n8774) );
  XNOR2_X1 U9837 ( .A(n8680), .B(n8681), .ZN(n8682) );
  OAI222_X1 U9838 ( .A1(n9637), .A2(n8809), .B1(n9635), .B2(n9307), .C1(n8682), 
        .C2(n9653), .ZN(n8775) );
  NAND2_X1 U9839 ( .A1(n8775), .A2(n10874), .ZN(n8685) );
  OAI22_X1 U9840 ( .A1(n10874), .A2(n5896), .B1(n9310), .B2(n9590), .ZN(n8683)
         );
  AOI21_X1 U9841 ( .B1(n9312), .B2(n10869), .A(n8683), .ZN(n8684) );
  OAI211_X1 U9842 ( .C1(n8774), .C2(n9629), .A(n8685), .B(n8684), .ZN(P2_U3217) );
  NOR2_X1 U9843 ( .A1(n8686), .A2(n9718), .ZN(n8688) );
  AOI211_X1 U9844 ( .C1(n9720), .C2(n8760), .A(n8688), .B(n8687), .ZN(n10987)
         );
  NAND2_X1 U9845 ( .A1(n9683), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8689) );
  OAI21_X1 U9846 ( .B1(n10987), .B2(n9683), .A(n8689), .ZN(P2_U3474) );
  NOR2_X1 U9847 ( .A1(n8690), .A2(n9718), .ZN(n8692) );
  AOI211_X1 U9848 ( .C1(n9720), .C2(n8706), .A(n8692), .B(n8691), .ZN(n10986)
         );
  OR2_X1 U9849 ( .A1(n10986), .A2(n9683), .ZN(n8693) );
  OAI21_X1 U9850 ( .B1(n9735), .B2(n8694), .A(n8693), .ZN(P2_U3473) );
  XOR2_X1 U9851 ( .A(n8695), .B(n8699), .Z(n8698) );
  OR2_X1 U9852 ( .A1(n9655), .A2(n9637), .ZN(n8697) );
  OR2_X1 U9853 ( .A1(n8809), .A2(n9635), .ZN(n8696) );
  AND2_X1 U9854 ( .A1(n8697), .A2(n8696), .ZN(n9362) );
  OAI21_X1 U9855 ( .B1(n8698), .B2(n9653), .A(n9362), .ZN(n9732) );
  INV_X1 U9856 ( .A(n9732), .ZN(n8705) );
  XNOR2_X1 U9857 ( .A(n8700), .B(n8699), .ZN(n9734) );
  INV_X1 U9858 ( .A(n8811), .ZN(n9780) );
  NOR2_X1 U9859 ( .A1(n9780), .A2(n9647), .ZN(n8703) );
  OAI22_X1 U9860 ( .A1(n10874), .A2(n8701), .B1(n9360), .B2(n9590), .ZN(n8702)
         );
  AOI211_X1 U9861 ( .C1(n9734), .C2(n9677), .A(n8703), .B(n8702), .ZN(n8704)
         );
  OAI21_X1 U9862 ( .B1(n8705), .B2(n9673), .A(n8704), .ZN(P2_U3215) );
  INV_X1 U9863 ( .A(n8706), .ZN(n8719) );
  XNOR2_X1 U9864 ( .A(n8706), .B(n7735), .ZN(n8758) );
  XNOR2_X1 U9865 ( .A(n8758), .B(n8767), .ZN(n8710) );
  OAI21_X1 U9866 ( .B1(n8710), .B2(n8709), .A(n8763), .ZN(n8711) );
  NAND2_X1 U9867 ( .A1(n8711), .A2(n5658), .ZN(n8718) );
  INV_X1 U9868 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8712) );
  OR2_X1 U9869 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8712), .ZN(n9452) );
  OAI21_X1 U9870 ( .B1(n9376), .B2(n8713), .A(n9452), .ZN(n8716) );
  NOR2_X1 U9871 ( .A1(n9377), .A2(n8714), .ZN(n8715) );
  AOI211_X1 U9872 ( .C1(n9380), .C2(n9391), .A(n8716), .B(n8715), .ZN(n8717)
         );
  OAI211_X1 U9873 ( .C1(n8719), .C2(n9383), .A(n8718), .B(n8717), .ZN(P2_U3155) );
  XNOR2_X1 U9874 ( .A(n8720), .B(n8725), .ZN(n8721) );
  OAI222_X1 U9875 ( .A1(n9635), .A2(n8806), .B1(n9637), .B2(n9316), .C1(n9653), 
        .C2(n8721), .ZN(n8730) );
  INV_X1 U9876 ( .A(n8722), .ZN(n8723) );
  AOI21_X1 U9877 ( .B1(n8725), .B2(n8724), .A(n8723), .ZN(n8734) );
  OAI22_X1 U9878 ( .A1(n8734), .A2(n9718), .B1(n8727), .B2(n8726), .ZN(n8728)
         );
  NOR2_X1 U9879 ( .A1(n8730), .A2(n8728), .ZN(n11016) );
  NAND2_X1 U9880 ( .A1(n9683), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8729) );
  OAI21_X1 U9881 ( .B1(n11016), .B2(n9683), .A(n8729), .ZN(P2_U3476) );
  NAND2_X1 U9882 ( .A1(n8730), .A2(n10874), .ZN(n8733) );
  OAI22_X1 U9883 ( .A1(n10874), .A2(n9501), .B1(n9319), .B2(n9590), .ZN(n8731)
         );
  AOI21_X1 U9884 ( .B1(n9321), .B2(n10869), .A(n8731), .ZN(n8732) );
  OAI211_X1 U9885 ( .C1(n8734), .C2(n9629), .A(n8733), .B(n8732), .ZN(P2_U3216) );
  NAND2_X1 U9886 ( .A1(n10957), .A2(n9948), .ZN(n8736) );
  OR2_X1 U9887 ( .A1(n10094), .A2(n7808), .ZN(n8735) );
  NAND2_X1 U9888 ( .A1(n8736), .A2(n8735), .ZN(n8737) );
  XNOR2_X1 U9889 ( .A(n8737), .B(n9899), .ZN(n9801) );
  NOR2_X1 U9890 ( .A1(n10094), .A2(n9901), .ZN(n8738) );
  AOI21_X1 U9891 ( .B1(n10957), .B2(n9863), .A(n8738), .ZN(n9800) );
  XNOR2_X1 U9892 ( .A(n9801), .B(n9800), .ZN(n8745) );
  INV_X1 U9893 ( .A(n9803), .ZN(n8743) );
  AOI21_X1 U9894 ( .B1(n8745), .B2(n8744), .A(n8743), .ZN(n8754) );
  INV_X1 U9895 ( .A(n10954), .ZN(n8751) );
  OR2_X1 U9896 ( .A1(n9924), .A2(n10462), .ZN(n8748) );
  OR2_X1 U9897 ( .A1(n8746), .A2(n10464), .ZN(n8747) );
  NAND2_X1 U9898 ( .A1(n8748), .A2(n8747), .ZN(n10944) );
  NAND2_X1 U9899 ( .A1(n10944), .A2(n10029), .ZN(n8750) );
  OAI211_X1 U9900 ( .C1(n10084), .C2(n8751), .A(n8750), .B(n8749), .ZN(n8752)
         );
  AOI21_X1 U9901 ( .B1(n10957), .B2(n10073), .A(n8752), .ZN(n8753) );
  OAI21_X1 U9902 ( .B1(n8754), .B2(n10064), .A(n8753), .ZN(P1_U3224) );
  INV_X1 U9903 ( .A(n8755), .ZN(n8782) );
  AOI21_X1 U9904 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n9790), .A(n8756), .ZN(
        n8757) );
  OAI21_X1 U9905 ( .B1(n8782), .B2(n9792), .A(n8757), .ZN(P2_U3268) );
  INV_X1 U9906 ( .A(n8760), .ZN(n8773) );
  INV_X1 U9907 ( .A(n8758), .ZN(n8759) );
  NAND2_X1 U9908 ( .A1(n8759), .A2(n8767), .ZN(n8761) );
  AND2_X1 U9909 ( .A1(n8763), .A2(n8761), .ZN(n8765) );
  XNOR2_X1 U9910 ( .A(n8760), .B(n7735), .ZN(n8803) );
  XNOR2_X1 U9911 ( .A(n8803), .B(n9307), .ZN(n8764) );
  NAND2_X1 U9912 ( .A1(n8763), .A2(n8762), .ZN(n8805) );
  OAI211_X1 U9913 ( .C1(n8765), .C2(n8764), .A(n5658), .B(n8805), .ZN(n8772)
         );
  OR2_X1 U9914 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8766), .ZN(n9470) );
  OAI21_X1 U9915 ( .B1(n9376), .B2(n8767), .A(n9470), .ZN(n8770) );
  NOR2_X1 U9916 ( .A1(n9377), .A2(n8768), .ZN(n8769) );
  AOI211_X1 U9917 ( .C1(n9380), .C2(n9390), .A(n8770), .B(n8769), .ZN(n8771)
         );
  OAI211_X1 U9918 ( .C1(n8773), .C2(n9383), .A(n8772), .B(n8771), .ZN(P2_U3181) );
  NOR2_X1 U9919 ( .A1(n8774), .A2(n9718), .ZN(n8776) );
  AOI211_X1 U9920 ( .C1(n9720), .C2(n9312), .A(n8776), .B(n8775), .ZN(n11014)
         );
  OR2_X1 U9921 ( .A1(n11014), .A2(n9683), .ZN(n8777) );
  OAI21_X1 U9922 ( .B1(n9735), .B2(n8778), .A(n8777), .ZN(P2_U3475) );
  INV_X1 U9923 ( .A(n8779), .ZN(n8781) );
  OAI222_X1 U9924 ( .A1(n8793), .A2(n9148), .B1(n8791), .B2(n8781), .C1(
        P1_U3086), .C2(n8780), .ZN(P1_U3329) );
  OAI222_X1 U9925 ( .A1(P2_U3151), .A2(n8784), .B1(n9792), .B2(n8781), .C1(
        n9783), .C2(n6061), .ZN(P2_U3269) );
  OAI222_X1 U9926 ( .A1(n8793), .A2(n9149), .B1(n8791), .B2(n8782), .C1(n7151), 
        .C2(P1_U3086), .ZN(P1_U3328) );
  AND2_X1 U9927 ( .A1(n8784), .A2(n8783), .ZN(n8785) );
  AOI22_X1 U9928 ( .A1(n8786), .A2(n5638), .B1(n8785), .B2(n6484), .ZN(
        P2_U3376) );
  INV_X1 U9929 ( .A(n8787), .ZN(n9793) );
  OAI222_X1 U9930 ( .A1(n8793), .A2(n10658), .B1(n8791), .B2(n9793), .C1(n8788), .C2(P1_U3086), .ZN(P1_U3327) );
  INV_X1 U9931 ( .A(n8789), .ZN(n9257) );
  OAI222_X1 U9932 ( .A1(n8793), .A2(n8792), .B1(n8791), .B2(n9257), .C1(n8790), 
        .C2(P1_U3086), .ZN(P1_U3326) );
  OAI21_X1 U9933 ( .B1(n8796), .B2(n8795), .A(n8794), .ZN(n8797) );
  NAND2_X1 U9934 ( .A1(n8797), .A2(n10081), .ZN(n8802) );
  OAI22_X1 U9935 ( .A1(n8799), .A2(n10464), .B1(n8798), .B2(n10462), .ZN(
        n10789) );
  AOI22_X1 U9936 ( .A1(n10789), .A2(n10029), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n8800), .ZN(n8801) );
  OAI211_X1 U9937 ( .C1(n7799), .C2(n10090), .A(n8802), .B(n8801), .ZN(
        P1_U3237) );
  INV_X1 U9938 ( .A(n8803), .ZN(n8804) );
  XNOR2_X1 U9939 ( .A(n9312), .B(n7766), .ZN(n8807) );
  NAND2_X1 U9940 ( .A1(n8807), .A2(n8806), .ZN(n9302) );
  NOR2_X1 U9941 ( .A1(n8807), .A2(n8806), .ZN(n9304) );
  XNOR2_X1 U9942 ( .A(n9321), .B(n7735), .ZN(n8808) );
  XNOR2_X1 U9943 ( .A(n8808), .B(n8809), .ZN(n9315) );
  INV_X1 U9944 ( .A(n8808), .ZN(n8810) );
  XNOR2_X1 U9945 ( .A(n8811), .B(n7735), .ZN(n8812) );
  XNOR2_X1 U9946 ( .A(n8812), .B(n9316), .ZN(n9358) );
  NAND2_X1 U9947 ( .A1(n8812), .A2(n9666), .ZN(n8813) );
  XNOR2_X1 U9948 ( .A(n9676), .B(n7766), .ZN(n9270) );
  INV_X1 U9949 ( .A(n9270), .ZN(n8814) );
  NAND2_X1 U9950 ( .A1(n8814), .A2(n9388), .ZN(n8815) );
  NAND2_X1 U9951 ( .A1(n9269), .A2(n8815), .ZN(n9339) );
  XNOR2_X1 U9952 ( .A(n9657), .B(n7735), .ZN(n8816) );
  XNOR2_X1 U9953 ( .A(n8816), .B(n9636), .ZN(n9338) );
  NAND2_X1 U9954 ( .A1(n9339), .A2(n9338), .ZN(n9337) );
  NAND2_X1 U9955 ( .A1(n8816), .A2(n9669), .ZN(n8817) );
  NAND2_X1 U9956 ( .A1(n9337), .A2(n8817), .ZN(n9288) );
  XNOR2_X1 U9957 ( .A(n9719), .B(n7735), .ZN(n8818) );
  XNOR2_X1 U9958 ( .A(n8818), .B(n9654), .ZN(n9287) );
  NAND2_X1 U9959 ( .A1(n8818), .A2(n5193), .ZN(n8819) );
  XNOR2_X1 U9960 ( .A(n8820), .B(n7735), .ZN(n8822) );
  XNOR2_X1 U9961 ( .A(n8822), .B(n9638), .ZN(n9348) );
  NAND2_X1 U9962 ( .A1(n8822), .A2(n9638), .ZN(n8823) );
  XNOR2_X1 U9963 ( .A(n9618), .B(n7766), .ZN(n8825) );
  INV_X1 U9964 ( .A(n8824), .ZN(n8826) );
  NAND2_X1 U9965 ( .A1(n8826), .A2(n8825), .ZN(n8827) );
  XNOR2_X1 U9966 ( .A(n9764), .B(n7735), .ZN(n8829) );
  XNOR2_X1 U9967 ( .A(n8829), .B(n9588), .ZN(n9326) );
  XNOR2_X1 U9968 ( .A(n9760), .B(n7735), .ZN(n9368) );
  NAND2_X1 U9969 ( .A1(n9325), .A2(n5708), .ZN(n8835) );
  NAND2_X1 U9970 ( .A1(n8829), .A2(n9588), .ZN(n9294) );
  INV_X1 U9971 ( .A(n9294), .ZN(n8833) );
  INV_X1 U9972 ( .A(n9368), .ZN(n8830) );
  AOI21_X1 U9973 ( .B1(n9387), .B2(n9294), .A(n8830), .ZN(n8832) );
  XNOR2_X1 U9974 ( .A(n9756), .B(n8831), .ZN(n8836) );
  XNOR2_X1 U9975 ( .A(n8836), .B(n9589), .ZN(n9371) );
  AOI211_X1 U9976 ( .C1(n9602), .C2(n8833), .A(n8832), .B(n9371), .ZN(n8834)
         );
  NAND2_X1 U9977 ( .A1(n8835), .A2(n8834), .ZN(n9372) );
  INV_X1 U9978 ( .A(n8836), .ZN(n8837) );
  XNOR2_X1 U9979 ( .A(n8841), .B(n7735), .ZN(n9278) );
  XNOR2_X1 U9980 ( .A(n9278), .B(n9576), .ZN(n9279) );
  NOR2_X1 U9981 ( .A1(n9377), .A2(n9568), .ZN(n8840) );
  AOI22_X1 U9982 ( .A1(n9330), .A2(n9386), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8838) );
  OAI21_X1 U9983 ( .B1(n10659), .B2(n9328), .A(n8838), .ZN(n8839) );
  AOI211_X1 U9984 ( .C1(n8841), .C2(n9353), .A(n8840), .B(n8839), .ZN(n8842)
         );
  XNOR2_X1 U9985 ( .A(n9044), .B(keyinput_3), .ZN(n8847) );
  XNOR2_X1 U9986 ( .A(n8843), .B(keyinput_2), .ZN(n8846) );
  XNOR2_X1 U9987 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_0), .ZN(n8845) );
  XNOR2_X1 U9988 ( .A(SI_31_), .B(keyinput_1), .ZN(n8844) );
  NOR4_X1 U9989 ( .A1(n8847), .A2(n8846), .A3(n8845), .A4(n8844), .ZN(n8854)
         );
  XNOR2_X1 U9990 ( .A(n9038), .B(keyinput_4), .ZN(n8851) );
  XNOR2_X1 U9991 ( .A(SI_26_), .B(keyinput_6), .ZN(n8850) );
  XNOR2_X1 U9992 ( .A(SI_27_), .B(keyinput_5), .ZN(n8849) );
  XNOR2_X1 U9993 ( .A(SI_25_), .B(keyinput_7), .ZN(n8848) );
  NAND4_X1 U9994 ( .A1(n8851), .A2(n8850), .A3(n8849), .A4(n8848), .ZN(n8853)
         );
  XNOR2_X1 U9995 ( .A(n9050), .B(keyinput_8), .ZN(n8852) );
  OAI21_X1 U9996 ( .B1(n8854), .B2(n8853), .A(n8852), .ZN(n8857) );
  XNOR2_X1 U9997 ( .A(n9055), .B(keyinput_10), .ZN(n8856) );
  XNOR2_X1 U9998 ( .A(n9054), .B(keyinput_9), .ZN(n8855) );
  NAND3_X1 U9999 ( .A1(n8857), .A2(n8856), .A3(n8855), .ZN(n8860) );
  XNOR2_X1 U10000 ( .A(SI_21_), .B(keyinput_11), .ZN(n8859) );
  XNOR2_X1 U10001 ( .A(SI_20_), .B(keyinput_12), .ZN(n8858) );
  NAND3_X1 U10002 ( .A1(n8860), .A2(n8859), .A3(n8858), .ZN(n8864) );
  XNOR2_X1 U10003 ( .A(SI_19_), .B(keyinput_13), .ZN(n8863) );
  XNOR2_X1 U10004 ( .A(n9064), .B(keyinput_15), .ZN(n8862) );
  XNOR2_X1 U10005 ( .A(SI_18_), .B(keyinput_14), .ZN(n8861) );
  AOI211_X1 U10006 ( .C1(n8864), .C2(n8863), .A(n8862), .B(n8861), .ZN(n8868)
         );
  XNOR2_X1 U10007 ( .A(SI_16_), .B(keyinput_16), .ZN(n8867) );
  XNOR2_X1 U10008 ( .A(SI_15_), .B(keyinput_17), .ZN(n8866) );
  XNOR2_X1 U10009 ( .A(SI_14_), .B(keyinput_18), .ZN(n8865) );
  OAI211_X1 U10010 ( .C1(n8868), .C2(n8867), .A(n8866), .B(n8865), .ZN(n8872)
         );
  XNOR2_X1 U10011 ( .A(SI_13_), .B(keyinput_19), .ZN(n8871) );
  XNOR2_X1 U10012 ( .A(n8869), .B(keyinput_20), .ZN(n8870) );
  AOI21_X1 U10013 ( .B1(n8872), .B2(n8871), .A(n8870), .ZN(n8876) );
  XNOR2_X1 U10014 ( .A(SI_11_), .B(keyinput_21), .ZN(n8875) );
  XNOR2_X1 U10015 ( .A(SI_9_), .B(keyinput_23), .ZN(n8874) );
  XNOR2_X1 U10016 ( .A(SI_10_), .B(keyinput_22), .ZN(n8873) );
  OAI211_X1 U10017 ( .C1(n8876), .C2(n8875), .A(n8874), .B(n8873), .ZN(n8888)
         );
  XOR2_X1 U10018 ( .A(SI_7_), .B(keyinput_25), .Z(n8882) );
  XNOR2_X1 U10019 ( .A(n8877), .B(keyinput_24), .ZN(n8881) );
  XNOR2_X1 U10020 ( .A(n8878), .B(keyinput_26), .ZN(n8880) );
  XNOR2_X1 U10021 ( .A(SI_5_), .B(keyinput_27), .ZN(n8879) );
  NOR4_X1 U10022 ( .A1(n8882), .A2(n8881), .A3(n8880), .A4(n8879), .ZN(n8887)
         );
  XNOR2_X1 U10023 ( .A(n8883), .B(keyinput_29), .ZN(n8886) );
  XNOR2_X1 U10024 ( .A(n8884), .B(keyinput_28), .ZN(n8885) );
  AOI211_X1 U10025 ( .C1(n8888), .C2(n8887), .A(n8886), .B(n8885), .ZN(n8891)
         );
  XNOR2_X1 U10026 ( .A(SI_2_), .B(keyinput_30), .ZN(n8890) );
  XOR2_X1 U10027 ( .A(SI_1_), .B(keyinput_31), .Z(n8889) );
  OAI21_X1 U10028 ( .B1(n8891), .B2(n8890), .A(n8889), .ZN(n8895) );
  XNOR2_X1 U10029 ( .A(P2_U3151), .B(keyinput_34), .ZN(n8894) );
  XNOR2_X1 U10030 ( .A(SI_0_), .B(keyinput_32), .ZN(n8893) );
  XNOR2_X1 U10031 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_33), .ZN(n8892) );
  NAND4_X1 U10032 ( .A1(n8895), .A2(n8894), .A3(n8893), .A4(n8892), .ZN(n8898)
         );
  XOR2_X1 U10033 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_35), .Z(n8897) );
  XOR2_X1 U10034 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_36), .Z(n8896) );
  AOI21_X1 U10035 ( .B1(n8898), .B2(n8897), .A(n8896), .ZN(n8905) );
  XOR2_X1 U10036 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_37), .Z(n8904) );
  XOR2_X1 U10037 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_40), .Z(n8902) );
  XOR2_X1 U10038 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_41), .Z(n8901) );
  XNOR2_X1 U10039 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_39), .ZN(n8900)
         );
  XNOR2_X1 U10040 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_38), .ZN(n8899)
         );
  NOR4_X1 U10041 ( .A1(n8902), .A2(n8901), .A3(n8900), .A4(n8899), .ZN(n8903)
         );
  OAI21_X1 U10042 ( .B1(n8905), .B2(n8904), .A(n8903), .ZN(n8908) );
  XNOR2_X1 U10043 ( .A(n9109), .B(keyinput_42), .ZN(n8907) );
  XNOR2_X1 U10044 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_43), .ZN(n8906) );
  NAND3_X1 U10045 ( .A1(n8908), .A2(n8907), .A3(n8906), .ZN(n8911) );
  XOR2_X1 U10046 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_44), .Z(n8910) );
  XNOR2_X1 U10047 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_45), .ZN(n8909)
         );
  AOI21_X1 U10048 ( .B1(n8911), .B2(n8910), .A(n8909), .ZN(n8918) );
  XOR2_X1 U10049 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_46), .Z(n8917) );
  XNOR2_X1 U10050 ( .A(n9116), .B(keyinput_49), .ZN(n8915) );
  XNOR2_X1 U10051 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_48), .ZN(n8914)
         );
  XNOR2_X1 U10052 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_50), .ZN(n8913)
         );
  XNOR2_X1 U10053 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput_47), .ZN(n8912)
         );
  NOR4_X1 U10054 ( .A1(n8915), .A2(n8914), .A3(n8913), .A4(n8912), .ZN(n8916)
         );
  OAI21_X1 U10055 ( .B1(n8918), .B2(n8917), .A(n8916), .ZN(n8921) );
  XNOR2_X1 U10056 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_51), .ZN(n8920)
         );
  XOR2_X1 U10057 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_52), .Z(n8919) );
  AOI21_X1 U10058 ( .B1(n8921), .B2(n8920), .A(n8919), .ZN(n8925) );
  XNOR2_X1 U10059 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput_53), .ZN(n8924) );
  XNOR2_X1 U10060 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .ZN(n8923) );
  XNOR2_X1 U10061 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_55), .ZN(n8922)
         );
  OAI211_X1 U10062 ( .C1(n8925), .C2(n8924), .A(n8923), .B(n8922), .ZN(n8928)
         );
  XOR2_X1 U10063 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_56), .Z(n8927) );
  XNOR2_X1 U10064 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_57), .ZN(n8926)
         );
  AOI21_X1 U10065 ( .B1(n8928), .B2(n8927), .A(n8926), .ZN(n8932) );
  XOR2_X1 U10066 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_58), .Z(n8931) );
  XNOR2_X1 U10067 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_60), .ZN(n8930)
         );
  XNOR2_X1 U10068 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_59), .ZN(n8929) );
  NOR4_X1 U10069 ( .A1(n8932), .A2(n8931), .A3(n8930), .A4(n8929), .ZN(n8936)
         );
  XNOR2_X1 U10070 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_61), .ZN(n8935) );
  XOR2_X1 U10071 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_62), .Z(n8934) );
  XNOR2_X1 U10072 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_63), .ZN(n8933)
         );
  OAI211_X1 U10073 ( .C1(n8936), .C2(n8935), .A(n8934), .B(n8933), .ZN(n8939)
         );
  XNOR2_X1 U10074 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_64), .ZN(n8938) );
  XNOR2_X1 U10075 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .ZN(n8937)
         );
  AOI21_X1 U10076 ( .B1(n8939), .B2(n8938), .A(n8937), .ZN(n8942) );
  XNOR2_X1 U10077 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_66), .ZN(n8941)
         );
  XNOR2_X1 U10078 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .ZN(n8940)
         );
  OAI21_X1 U10079 ( .B1(n8942), .B2(n8941), .A(n8940), .ZN(n8946) );
  XOR2_X1 U10080 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .Z(n8945) );
  XNOR2_X1 U10081 ( .A(n9149), .B(keyinput_69), .ZN(n8944) );
  XNOR2_X1 U10082 ( .A(n9148), .B(keyinput_70), .ZN(n8943) );
  AOI211_X1 U10083 ( .C1(n8946), .C2(n8945), .A(n8944), .B(n8943), .ZN(n8954)
         );
  XNOR2_X1 U10084 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .ZN(n8953)
         );
  XNOR2_X1 U10085 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .ZN(n8952)
         );
  XOR2_X1 U10086 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .Z(n8950) );
  XNOR2_X1 U10087 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .ZN(n8949)
         );
  XNOR2_X1 U10088 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_76), .ZN(n8948)
         );
  XNOR2_X1 U10089 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .ZN(n8947)
         );
  NAND4_X1 U10090 ( .A1(n8950), .A2(n8949), .A3(n8948), .A4(n8947), .ZN(n8951)
         );
  NOR4_X1 U10091 ( .A1(n8954), .A2(n8953), .A3(n8952), .A4(n8951), .ZN(n8957)
         );
  XNOR2_X1 U10092 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .ZN(n8956)
         );
  XOR2_X1 U10093 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .Z(n8955) );
  OAI21_X1 U10094 ( .B1(n8957), .B2(n8956), .A(n8955), .ZN(n8963) );
  XOR2_X1 U10095 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .Z(n8961) );
  XNOR2_X1 U10096 ( .A(n9168), .B(keyinput_79), .ZN(n8960) );
  XNOR2_X1 U10097 ( .A(n9169), .B(keyinput_80), .ZN(n8959) );
  XNOR2_X1 U10098 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_82), .ZN(n8958)
         );
  NOR4_X1 U10099 ( .A1(n8961), .A2(n8960), .A3(n8959), .A4(n8958), .ZN(n8962)
         );
  NAND2_X1 U10100 ( .A1(n8963), .A2(n8962), .ZN(n8970) );
  INV_X1 U10101 ( .A(keyinput_84), .ZN(n8964) );
  XNOR2_X1 U10102 ( .A(n8964), .B(P2_DATAO_REG_12__SCAN_IN), .ZN(n8969) );
  OAI22_X1 U10103 ( .A1(n8966), .A2(keyinput_83), .B1(keyinput_85), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n8965) );
  AOI21_X1 U10104 ( .B1(n8966), .B2(keyinput_83), .A(n8965), .ZN(n8968) );
  NAND2_X1 U10105 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput_85), .ZN(n8967) );
  NAND4_X1 U10106 ( .A1(n8970), .A2(n8969), .A3(n8968), .A4(n8967), .ZN(n8973)
         );
  XOR2_X1 U10107 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_86), .Z(n8972) );
  XNOR2_X1 U10108 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_87), .ZN(n8971)
         );
  AOI21_X1 U10109 ( .B1(n8973), .B2(n8972), .A(n8971), .ZN(n8977) );
  XOR2_X1 U10110 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_90), .Z(n8976) );
  XNOR2_X1 U10111 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .ZN(n8975)
         );
  XNOR2_X1 U10112 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .ZN(n8974)
         );
  NOR4_X1 U10113 ( .A1(n8977), .A2(n8976), .A3(n8975), .A4(n8974), .ZN(n8980)
         );
  XNOR2_X1 U10114 ( .A(n9189), .B(keyinput_92), .ZN(n8979) );
  XNOR2_X1 U10115 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_91), .ZN(n8978) );
  NOR3_X1 U10116 ( .A1(n8980), .A2(n8979), .A3(n8978), .ZN(n8983) );
  XOR2_X1 U10117 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_93), .Z(n8982) );
  XOR2_X1 U10118 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_94), .Z(n8981) );
  NOR3_X1 U10119 ( .A1(n8983), .A2(n8982), .A3(n8981), .ZN(n8993) );
  INV_X1 U10120 ( .A(keyinput_97), .ZN(n8989) );
  INV_X1 U10121 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8988) );
  XNOR2_X1 U10122 ( .A(n8984), .B(keyinput_96), .ZN(n8987) );
  INV_X1 U10123 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9197) );
  OAI22_X1 U10124 ( .A1(n9197), .A2(keyinput_95), .B1(keyinput_97), .B2(
        P1_IR_REG_7__SCAN_IN), .ZN(n8985) );
  AOI21_X1 U10125 ( .B1(n9197), .B2(keyinput_95), .A(n8985), .ZN(n8986) );
  OAI211_X1 U10126 ( .C1(n8989), .C2(n8988), .A(n8987), .B(n8986), .ZN(n8992)
         );
  XOR2_X1 U10127 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_98), .Z(n8991) );
  XNOR2_X1 U10128 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_99), .ZN(n8990) );
  OAI211_X1 U10129 ( .C1(n8993), .C2(n8992), .A(n8991), .B(n8990), .ZN(n9000)
         );
  XNOR2_X1 U10130 ( .A(n8994), .B(keyinput_101), .ZN(n8996) );
  XNOR2_X1 U10131 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_100), .ZN(n8995) );
  NOR2_X1 U10132 ( .A1(n8996), .A2(n8995), .ZN(n8999) );
  XNOR2_X1 U10133 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_103), .ZN(n8998) );
  XNOR2_X1 U10134 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_102), .ZN(n8997) );
  AOI211_X1 U10135 ( .C1(n9000), .C2(n8999), .A(n8998), .B(n8997), .ZN(n9005)
         );
  XNOR2_X1 U10136 ( .A(n9001), .B(keyinput_104), .ZN(n9004) );
  XNOR2_X1 U10137 ( .A(n9211), .B(keyinput_106), .ZN(n9003) );
  XNOR2_X1 U10138 ( .A(n9212), .B(keyinput_105), .ZN(n9002) );
  OAI211_X1 U10139 ( .C1(n9005), .C2(n9004), .A(n9003), .B(n9002), .ZN(n9008)
         );
  XNOR2_X1 U10140 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_107), .ZN(n9007) );
  XNOR2_X1 U10141 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_108), .ZN(n9006) );
  NAND3_X1 U10142 ( .A1(n9008), .A2(n9007), .A3(n9006), .ZN(n9016) );
  XNOR2_X1 U10143 ( .A(n9009), .B(keyinput_112), .ZN(n9013) );
  XNOR2_X1 U10144 ( .A(n9221), .B(keyinput_111), .ZN(n9012) );
  XNOR2_X1 U10145 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_109), .ZN(n9011) );
  XNOR2_X1 U10146 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_110), .ZN(n9010) );
  NOR4_X1 U10147 ( .A1(n9013), .A2(n9012), .A3(n9011), .A4(n9010), .ZN(n9015)
         );
  XNOR2_X1 U10148 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_113), .ZN(n9014) );
  AOI21_X1 U10149 ( .B1(n9016), .B2(n9015), .A(n9014), .ZN(n9020) );
  XNOR2_X1 U10150 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_114), .ZN(n9019) );
  XNOR2_X1 U10151 ( .A(n9017), .B(keyinput_115), .ZN(n9018) );
  OAI21_X1 U10152 ( .B1(n9020), .B2(n9019), .A(n9018), .ZN(n9024) );
  XNOR2_X1 U10153 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_116), .ZN(n9023) );
  XNOR2_X1 U10154 ( .A(n9021), .B(keyinput_117), .ZN(n9022) );
  AOI21_X1 U10155 ( .B1(n9024), .B2(n9023), .A(n9022), .ZN(n9028) );
  XNOR2_X1 U10156 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_118), .ZN(n9027) );
  XNOR2_X1 U10157 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_119), .ZN(n9026) );
  XNOR2_X1 U10158 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_120), .ZN(n9025) );
  OAI211_X1 U10159 ( .C1(n9028), .C2(n9027), .A(n9026), .B(n9025), .ZN(n9036)
         );
  XOR2_X1 U10160 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_123), .Z(n9032) );
  XOR2_X1 U10161 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_121), .Z(n9031) );
  XNOR2_X1 U10162 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_122), .ZN(n9030) );
  XNOR2_X1 U10163 ( .A(P1_D_REG_2__SCAN_IN), .B(keyinput_124), .ZN(n9029) );
  NOR4_X1 U10164 ( .A1(n9032), .A2(n9031), .A3(n9030), .A4(n9029), .ZN(n9035)
         );
  INV_X1 U10165 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10588) );
  XNOR2_X1 U10166 ( .A(n10588), .B(keyinput_126), .ZN(n9034) );
  XNOR2_X1 U10167 ( .A(P1_D_REG_3__SCAN_IN), .B(keyinput_125), .ZN(n9033) );
  AOI211_X1 U10168 ( .C1(n9036), .C2(n9035), .A(n9034), .B(n9033), .ZN(n9253)
         );
  XNOR2_X1 U10169 ( .A(keyinput_255), .B(keyinput_127), .ZN(n9252) );
  XOR2_X1 U10170 ( .A(keyinput_255), .B(P1_D_REG_5__SCAN_IN), .Z(n9251) );
  XNOR2_X1 U10171 ( .A(n9037), .B(keyinput_134), .ZN(n9043) );
  XNOR2_X1 U10172 ( .A(n9038), .B(keyinput_132), .ZN(n9042) );
  XNOR2_X1 U10173 ( .A(n9039), .B(keyinput_133), .ZN(n9041) );
  XNOR2_X1 U10174 ( .A(SI_25_), .B(keyinput_135), .ZN(n9040) );
  NOR4_X1 U10175 ( .A1(n9043), .A2(n9042), .A3(n9041), .A4(n9040), .ZN(n9053)
         );
  XOR2_X1 U10176 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_128), .Z(n9049) );
  XNOR2_X1 U10177 ( .A(n9044), .B(keyinput_131), .ZN(n9048) );
  XNOR2_X1 U10178 ( .A(n9045), .B(keyinput_129), .ZN(n9047) );
  XNOR2_X1 U10179 ( .A(SI_30_), .B(keyinput_130), .ZN(n9046) );
  NAND4_X1 U10180 ( .A1(n9049), .A2(n9048), .A3(n9047), .A4(n9046), .ZN(n9052)
         );
  XNOR2_X1 U10181 ( .A(n9050), .B(keyinput_136), .ZN(n9051) );
  AOI21_X1 U10182 ( .B1(n9053), .B2(n9052), .A(n9051), .ZN(n9058) );
  XNOR2_X1 U10183 ( .A(n9054), .B(keyinput_137), .ZN(n9057) );
  XNOR2_X1 U10184 ( .A(n9055), .B(keyinput_138), .ZN(n9056) );
  NOR3_X1 U10185 ( .A1(n9058), .A2(n9057), .A3(n9056), .ZN(n9063) );
  XNOR2_X1 U10186 ( .A(n9059), .B(keyinput_139), .ZN(n9062) );
  XNOR2_X1 U10187 ( .A(n9060), .B(keyinput_140), .ZN(n9061) );
  NOR3_X1 U10188 ( .A1(n9063), .A2(n9062), .A3(n9061), .ZN(n9068) );
  XNOR2_X1 U10189 ( .A(SI_19_), .B(keyinput_141), .ZN(n9067) );
  XNOR2_X1 U10190 ( .A(n9064), .B(keyinput_143), .ZN(n9066) );
  XNOR2_X1 U10191 ( .A(SI_18_), .B(keyinput_142), .ZN(n9065) );
  OAI211_X1 U10192 ( .C1(n9068), .C2(n9067), .A(n9066), .B(n9065), .ZN(n9073)
         );
  XNOR2_X1 U10193 ( .A(SI_16_), .B(keyinput_144), .ZN(n9072) );
  XNOR2_X1 U10194 ( .A(n9069), .B(keyinput_146), .ZN(n9071) );
  XNOR2_X1 U10195 ( .A(SI_15_), .B(keyinput_145), .ZN(n9070) );
  AOI211_X1 U10196 ( .C1(n9073), .C2(n9072), .A(n9071), .B(n9070), .ZN(n9076)
         );
  XNOR2_X1 U10197 ( .A(SI_13_), .B(keyinput_147), .ZN(n9075) );
  XNOR2_X1 U10198 ( .A(SI_12_), .B(keyinput_148), .ZN(n9074) );
  OAI21_X1 U10199 ( .B1(n9076), .B2(n9075), .A(n9074), .ZN(n9082) );
  XNOR2_X1 U10200 ( .A(SI_11_), .B(keyinput_149), .ZN(n9081) );
  XNOR2_X1 U10201 ( .A(n9077), .B(keyinput_151), .ZN(n9080) );
  XNOR2_X1 U10202 ( .A(n9078), .B(keyinput_150), .ZN(n9079) );
  AOI211_X1 U10203 ( .C1(n9082), .C2(n9081), .A(n9080), .B(n9079), .ZN(n9091)
         );
  XNOR2_X1 U10204 ( .A(n9083), .B(keyinput_155), .ZN(n9087) );
  XNOR2_X1 U10205 ( .A(SI_7_), .B(keyinput_153), .ZN(n9086) );
  XNOR2_X1 U10206 ( .A(SI_8_), .B(keyinput_152), .ZN(n9085) );
  XNOR2_X1 U10207 ( .A(SI_6_), .B(keyinput_154), .ZN(n9084) );
  NAND4_X1 U10208 ( .A1(n9087), .A2(n9086), .A3(n9085), .A4(n9084), .ZN(n9090)
         );
  XNOR2_X1 U10209 ( .A(SI_3_), .B(keyinput_157), .ZN(n9089) );
  XNOR2_X1 U10210 ( .A(SI_4_), .B(keyinput_156), .ZN(n9088) );
  OAI211_X1 U10211 ( .C1(n9091), .C2(n9090), .A(n9089), .B(n9088), .ZN(n9094)
         );
  XNOR2_X1 U10212 ( .A(SI_2_), .B(keyinput_158), .ZN(n9093) );
  XNOR2_X1 U10213 ( .A(SI_1_), .B(keyinput_159), .ZN(n9092) );
  AOI21_X1 U10214 ( .B1(n9094), .B2(n9093), .A(n9092), .ZN(n9098) );
  XNOR2_X1 U10215 ( .A(P2_U3151), .B(keyinput_162), .ZN(n9097) );
  XOR2_X1 U10216 ( .A(SI_0_), .B(keyinput_160), .Z(n9096) );
  XNOR2_X1 U10217 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_161), .ZN(n9095) );
  NOR4_X1 U10218 ( .A1(n9098), .A2(n9097), .A3(n9096), .A4(n9095), .ZN(n9101)
         );
  XNOR2_X1 U10219 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_163), .ZN(n9100)
         );
  XNOR2_X1 U10220 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_164), .ZN(n9099)
         );
  OAI21_X1 U10221 ( .B1(n9101), .B2(n9100), .A(n9099), .ZN(n9108) );
  XOR2_X1 U10222 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_165), .Z(n9107) );
  XOR2_X1 U10223 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_168), .Z(n9105) );
  XOR2_X1 U10224 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_166), .Z(n9104) );
  XNOR2_X1 U10225 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_167), .ZN(n9103)
         );
  XNOR2_X1 U10226 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_169), .ZN(n9102)
         );
  NAND4_X1 U10227 ( .A1(n9105), .A2(n9104), .A3(n9103), .A4(n9102), .ZN(n9106)
         );
  AOI21_X1 U10228 ( .B1(n9108), .B2(n9107), .A(n9106), .ZN(n9112) );
  XNOR2_X1 U10229 ( .A(n9109), .B(keyinput_170), .ZN(n9111) );
  XNOR2_X1 U10230 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_171), .ZN(n9110)
         );
  NOR3_X1 U10231 ( .A1(n9112), .A2(n9111), .A3(n9110), .ZN(n9115) );
  XOR2_X1 U10232 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_172), .Z(n9114) );
  XNOR2_X1 U10233 ( .A(n9289), .B(keyinput_173), .ZN(n9113) );
  OAI21_X1 U10234 ( .B1(n9115), .B2(n9114), .A(n9113), .ZN(n9123) );
  XNOR2_X1 U10235 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_174), .ZN(n9122)
         );
  XOR2_X1 U10236 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_176), .Z(n9120) );
  XNOR2_X1 U10237 ( .A(n9116), .B(keyinput_177), .ZN(n9119) );
  XNOR2_X1 U10238 ( .A(n9296), .B(keyinput_175), .ZN(n9118) );
  XNOR2_X1 U10239 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_178), .ZN(n9117)
         );
  NAND4_X1 U10240 ( .A1(n9120), .A2(n9119), .A3(n9118), .A4(n9117), .ZN(n9121)
         );
  AOI21_X1 U10241 ( .B1(n9123), .B2(n9122), .A(n9121), .ZN(n9126) );
  XNOR2_X1 U10242 ( .A(n9327), .B(keyinput_179), .ZN(n9125) );
  XNOR2_X1 U10243 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_180), .ZN(n9124)
         );
  OAI21_X1 U10244 ( .B1(n9126), .B2(n9125), .A(n9124), .ZN(n9130) );
  XNOR2_X1 U10245 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput_181), .ZN(n9129)
         );
  XOR2_X1 U10246 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_183), .Z(n9128) );
  XNOR2_X1 U10247 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_182), .ZN(n9127)
         );
  AOI211_X1 U10248 ( .C1(n9130), .C2(n9129), .A(n9128), .B(n9127), .ZN(n9133)
         );
  XOR2_X1 U10249 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_184), .Z(n9132) );
  XOR2_X1 U10250 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_185), .Z(n9131) );
  OAI21_X1 U10251 ( .B1(n9133), .B2(n9132), .A(n9131), .ZN(n9137) );
  XOR2_X1 U10252 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_187), .Z(n9136) );
  XOR2_X1 U10253 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_186), .Z(n9135) );
  XNOR2_X1 U10254 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_188), .ZN(n9134)
         );
  NAND4_X1 U10255 ( .A1(n9137), .A2(n9136), .A3(n9135), .A4(n9134), .ZN(n9141)
         );
  XNOR2_X1 U10256 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_189), .ZN(n9140)
         );
  XOR2_X1 U10257 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_191), .Z(n9139) );
  XNOR2_X1 U10258 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_190), .ZN(n9138)
         );
  AOI211_X1 U10259 ( .C1(n9141), .C2(n9140), .A(n9139), .B(n9138), .ZN(n9144)
         );
  XOR2_X1 U10260 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_192), .Z(n9143) );
  XOR2_X1 U10261 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_193), .Z(n9142)
         );
  OAI21_X1 U10262 ( .B1(n9144), .B2(n9143), .A(n9142), .ZN(n9147) );
  XNOR2_X1 U10263 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_194), .ZN(n9146)
         );
  XNOR2_X1 U10264 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_195), .ZN(n9145)
         );
  AOI21_X1 U10265 ( .B1(n9147), .B2(n9146), .A(n9145), .ZN(n9153) );
  XNOR2_X1 U10266 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_196), .ZN(n9152)
         );
  XNOR2_X1 U10267 ( .A(n9148), .B(keyinput_198), .ZN(n9151) );
  XNOR2_X1 U10268 ( .A(n9149), .B(keyinput_197), .ZN(n9150) );
  OAI211_X1 U10269 ( .C1(n9153), .C2(n9152), .A(n9151), .B(n9150), .ZN(n9164)
         );
  XOR2_X1 U10270 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_203), .Z(n9163)
         );
  XNOR2_X1 U10271 ( .A(n9154), .B(keyinput_200), .ZN(n9162) );
  XNOR2_X1 U10272 ( .A(n9155), .B(keyinput_201), .ZN(n9160) );
  XNOR2_X1 U10273 ( .A(n9156), .B(keyinput_202), .ZN(n9159) );
  XOR2_X1 U10274 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_199), .Z(n9158)
         );
  XNOR2_X1 U10275 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_204), .ZN(n9157)
         );
  NOR4_X1 U10276 ( .A1(n9160), .A2(n9159), .A3(n9158), .A4(n9157), .ZN(n9161)
         );
  NAND4_X1 U10277 ( .A1(n9164), .A2(n9163), .A3(n9162), .A4(n9161), .ZN(n9167)
         );
  XNOR2_X1 U10278 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_205), .ZN(n9166)
         );
  XNOR2_X1 U10279 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_206), .ZN(n9165)
         );
  AOI21_X1 U10280 ( .B1(n9167), .B2(n9166), .A(n9165), .ZN(n9179) );
  XOR2_X1 U10281 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_209), .Z(n9173)
         );
  XNOR2_X1 U10282 ( .A(n9168), .B(keyinput_207), .ZN(n9172) );
  XNOR2_X1 U10283 ( .A(n9169), .B(keyinput_208), .ZN(n9171) );
  XNOR2_X1 U10284 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_210), .ZN(n9170)
         );
  NAND4_X1 U10285 ( .A1(n9173), .A2(n9172), .A3(n9171), .A4(n9170), .ZN(n9178)
         );
  XOR2_X1 U10286 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_211), .Z(n9176)
         );
  XNOR2_X1 U10287 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_212), .ZN(n9175)
         );
  XNOR2_X1 U10288 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_213), .ZN(n9174)
         );
  NOR3_X1 U10289 ( .A1(n9176), .A2(n9175), .A3(n9174), .ZN(n9177) );
  OAI21_X1 U10290 ( .B1(n9179), .B2(n9178), .A(n9177), .ZN(n9183) );
  XOR2_X1 U10291 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_214), .Z(n9182)
         );
  XNOR2_X1 U10292 ( .A(n9180), .B(keyinput_215), .ZN(n9181) );
  AOI21_X1 U10293 ( .B1(n9183), .B2(n9182), .A(n9181), .ZN(n9193) );
  INV_X1 U10294 ( .A(keyinput_217), .ZN(n9188) );
  XOR2_X1 U10295 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_218), .Z(n9186) );
  OAI22_X1 U10296 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput_216), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_217), .ZN(n9184) );
  AOI21_X1 U10297 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_216), .A(n9184), 
        .ZN(n9185) );
  OAI211_X1 U10298 ( .C1(n9188), .C2(n9187), .A(n9186), .B(n9185), .ZN(n9192)
         );
  XOR2_X1 U10299 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_219), .Z(n9191) );
  XNOR2_X1 U10300 ( .A(n9189), .B(keyinput_220), .ZN(n9190) );
  OAI211_X1 U10301 ( .C1(n9193), .C2(n9192), .A(n9191), .B(n9190), .ZN(n9196)
         );
  XOR2_X1 U10302 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_222), .Z(n9195) );
  XNOR2_X1 U10303 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_221), .ZN(n9194) );
  NAND3_X1 U10304 ( .A1(n9196), .A2(n9195), .A3(n9194), .ZN(n9201) );
  XNOR2_X1 U10305 ( .A(n9197), .B(keyinput_223), .ZN(n9200) );
  XOR2_X1 U10306 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_225), .Z(n9199) );
  XNOR2_X1 U10307 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_224), .ZN(n9198) );
  NAND4_X1 U10308 ( .A1(n9201), .A2(n9200), .A3(n9199), .A4(n9198), .ZN(n9204)
         );
  XNOR2_X1 U10309 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_226), .ZN(n9203) );
  XNOR2_X1 U10310 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_227), .ZN(n9202) );
  NAND3_X1 U10311 ( .A1(n9204), .A2(n9203), .A3(n9202), .ZN(n9207) );
  XNOR2_X1 U10312 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_229), .ZN(n9206) );
  XNOR2_X1 U10313 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_228), .ZN(n9205) );
  NAND3_X1 U10314 ( .A1(n9207), .A2(n9206), .A3(n9205), .ZN(n9210) );
  XOR2_X1 U10315 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_230), .Z(n9209) );
  XNOR2_X1 U10316 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_231), .ZN(n9208) );
  NAND3_X1 U10317 ( .A1(n9210), .A2(n9209), .A3(n9208), .ZN(n9216) );
  XNOR2_X1 U10318 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_232), .ZN(n9215) );
  XNOR2_X1 U10319 ( .A(n9211), .B(keyinput_234), .ZN(n9214) );
  XNOR2_X1 U10320 ( .A(n9212), .B(keyinput_233), .ZN(n9213) );
  AOI211_X1 U10321 ( .C1(n9216), .C2(n9215), .A(n9214), .B(n9213), .ZN(n9220)
         );
  XNOR2_X1 U10322 ( .A(n9217), .B(keyinput_235), .ZN(n9219) );
  XNOR2_X1 U10323 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_236), .ZN(n9218) );
  NOR3_X1 U10324 ( .A1(n9220), .A2(n9219), .A3(n9218), .ZN(n9229) );
  XNOR2_X1 U10325 ( .A(n9221), .B(keyinput_239), .ZN(n9225) );
  XNOR2_X1 U10326 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_240), .ZN(n9224) );
  XNOR2_X1 U10327 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_237), .ZN(n9223) );
  XNOR2_X1 U10328 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_238), .ZN(n9222) );
  NAND4_X1 U10329 ( .A1(n9225), .A2(n9224), .A3(n9223), .A4(n9222), .ZN(n9228)
         );
  XNOR2_X1 U10330 ( .A(n9226), .B(keyinput_241), .ZN(n9227) );
  OAI21_X1 U10331 ( .B1(n9229), .B2(n9228), .A(n9227), .ZN(n9232) );
  XOR2_X1 U10332 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_242), .Z(n9231) );
  XNOR2_X1 U10333 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_243), .ZN(n9230) );
  AOI21_X1 U10334 ( .B1(n9232), .B2(n9231), .A(n9230), .ZN(n9235) );
  XOR2_X1 U10335 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_244), .Z(n9234) );
  XNOR2_X1 U10336 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_245), .ZN(n9233) );
  OAI21_X1 U10337 ( .B1(n9235), .B2(n9234), .A(n9233), .ZN(n9241) );
  XNOR2_X1 U10338 ( .A(n9236), .B(keyinput_246), .ZN(n9240) );
  XNOR2_X1 U10339 ( .A(n9237), .B(keyinput_247), .ZN(n9239) );
  XNOR2_X1 U10340 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_248), .ZN(n9238) );
  AOI211_X1 U10341 ( .C1(n9241), .C2(n9240), .A(n9239), .B(n9238), .ZN(n9249)
         );
  XOR2_X1 U10342 ( .A(P1_D_REG_2__SCAN_IN), .B(keyinput_252), .Z(n9245) );
  XOR2_X1 U10343 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_250), .Z(n9244) );
  XOR2_X1 U10344 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_251), .Z(n9243) );
  XNOR2_X1 U10345 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_249), .ZN(n9242) );
  NAND4_X1 U10346 ( .A1(n9245), .A2(n9244), .A3(n9243), .A4(n9242), .ZN(n9248)
         );
  XOR2_X1 U10347 ( .A(P1_D_REG_3__SCAN_IN), .B(keyinput_253), .Z(n9247) );
  XNOR2_X1 U10348 ( .A(P1_D_REG_4__SCAN_IN), .B(keyinput_254), .ZN(n9246) );
  OAI211_X1 U10349 ( .C1(n9249), .C2(n9248), .A(n9247), .B(n9246), .ZN(n9250)
         );
  OAI211_X1 U10350 ( .C1(n9253), .C2(n9252), .A(n9251), .B(n9250), .ZN(n9254)
         );
  OAI222_X1 U10351 ( .A1(n9792), .A2(n9257), .B1(n9256), .B2(P2_U3151), .C1(
        n9255), .C2(n9783), .ZN(P2_U3266) );
  INV_X1 U10352 ( .A(n9258), .ZN(n10586) );
  OAI222_X1 U10353 ( .A1(n9261), .A2(n9260), .B1(n9792), .B2(n10586), .C1(
        P2_U3151), .C2(n9259), .ZN(P2_U3265) );
  OAI211_X1 U10354 ( .C1(n9263), .C2(n9622), .A(n9262), .B(n5658), .ZN(n9268)
         );
  INV_X1 U10355 ( .A(n9264), .ZN(n9616) );
  AOI22_X1 U10356 ( .A1(n9380), .A2(n9612), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n9265) );
  OAI21_X1 U10357 ( .B1(n9638), .B2(n9376), .A(n9265), .ZN(n9266) );
  AOI21_X1 U10358 ( .B1(n9616), .B2(n9364), .A(n9266), .ZN(n9267) );
  OAI211_X1 U10359 ( .C1(n9618), .C2(n9383), .A(n9268), .B(n9267), .ZN(
        P2_U3156) );
  INV_X1 U10360 ( .A(n9674), .ZN(n9775) );
  OAI211_X1 U10361 ( .C1(n9271), .C2(n9270), .A(n9269), .B(n5658), .ZN(n9277)
         );
  INV_X1 U10362 ( .A(n9272), .ZN(n9672) );
  NAND2_X1 U10363 ( .A1(n9330), .A2(n9666), .ZN(n9274) );
  OAI211_X1 U10364 ( .C1(n9328), .C2(n9636), .A(n9274), .B(n9273), .ZN(n9275)
         );
  AOI21_X1 U10365 ( .B1(n9672), .B2(n9364), .A(n9275), .ZN(n9276) );
  OAI211_X1 U10366 ( .C1(n9775), .C2(n9383), .A(n9277), .B(n9276), .ZN(
        P2_U3159) );
  XNOR2_X1 U10367 ( .A(n9556), .B(n7735), .ZN(n9280) );
  INV_X1 U10368 ( .A(n9281), .ZN(n9554) );
  NAND2_X1 U10369 ( .A1(n9364), .A2(n9554), .ZN(n9283) );
  AOI22_X1 U10370 ( .A1(n9330), .A2(n9385), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n9282) );
  OAI211_X1 U10371 ( .C1(n9550), .C2(n9328), .A(n9283), .B(n9282), .ZN(n9284)
         );
  AOI21_X1 U10372 ( .B1(n9555), .B2(n9353), .A(n9284), .ZN(n9285) );
  OAI211_X1 U10373 ( .C1(n9288), .C2(n9287), .A(n9286), .B(n5658), .ZN(n9293)
         );
  OAI22_X1 U10374 ( .A1(n9328), .A2(n9638), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9289), .ZN(n9291) );
  NOR2_X1 U10375 ( .A1(n9376), .A2(n9636), .ZN(n9290) );
  AOI211_X1 U10376 ( .C1(n9645), .C2(n9364), .A(n9291), .B(n9290), .ZN(n9292)
         );
  OAI211_X1 U10377 ( .C1(n9648), .C2(n9383), .A(n9293), .B(n9292), .ZN(
        P2_U3163) );
  XNOR2_X1 U10378 ( .A(n9368), .B(n9387), .ZN(n9369) );
  NAND2_X1 U10379 ( .A1(n9295), .A2(n9294), .ZN(n9370) );
  XOR2_X1 U10380 ( .A(n9369), .B(n9370), .Z(n9301) );
  OAI22_X1 U10381 ( .A1(n9328), .A2(n9589), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9296), .ZN(n9297) );
  AOI21_X1 U10382 ( .B1(n9330), .B2(n9612), .A(n9297), .ZN(n9298) );
  OAI21_X1 U10383 ( .B1(n9377), .B2(n9591), .A(n9298), .ZN(n9299) );
  AOI21_X1 U10384 ( .B1(n6393), .B2(n9353), .A(n9299), .ZN(n9300) );
  OAI21_X1 U10385 ( .B1(n9301), .B2(n9355), .A(n9300), .ZN(P2_U3165) );
  INV_X1 U10386 ( .A(n9302), .ZN(n9303) );
  NOR2_X1 U10387 ( .A1(n9304), .A2(n9303), .ZN(n9305) );
  XNOR2_X1 U10388 ( .A(n9306), .B(n9305), .ZN(n9314) );
  NAND2_X1 U10389 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9486) );
  OAI21_X1 U10390 ( .B1(n9376), .B2(n9307), .A(n9486), .ZN(n9308) );
  AOI21_X1 U10391 ( .B1(n9380), .B2(n9389), .A(n9308), .ZN(n9309) );
  OAI21_X1 U10392 ( .B1(n9310), .B2(n9377), .A(n9309), .ZN(n9311) );
  AOI21_X1 U10393 ( .B1(n9312), .B2(n9353), .A(n9311), .ZN(n9313) );
  OAI21_X1 U10394 ( .B1(n9314), .B2(n9355), .A(n9313), .ZN(P2_U3166) );
  XOR2_X1 U10395 ( .A(n9315), .B(n5177), .Z(n9323) );
  NAND2_X1 U10396 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9502) );
  OAI21_X1 U10397 ( .B1(n9328), .B2(n9316), .A(n9502), .ZN(n9317) );
  AOI21_X1 U10398 ( .B1(n9330), .B2(n9390), .A(n9317), .ZN(n9318) );
  OAI21_X1 U10399 ( .B1(n9377), .B2(n9319), .A(n9318), .ZN(n9320) );
  AOI21_X1 U10400 ( .B1(n9321), .B2(n9353), .A(n9320), .ZN(n9322) );
  OAI21_X1 U10401 ( .B1(n9323), .B2(n9355), .A(n9322), .ZN(P2_U3168) );
  AOI21_X1 U10402 ( .B1(n9326), .B2(n9324), .A(n9325), .ZN(n9336) );
  OAI22_X1 U10403 ( .A1(n9328), .A2(n9602), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9327), .ZN(n9329) );
  AOI21_X1 U10404 ( .B1(n9330), .B2(n9622), .A(n9329), .ZN(n9331) );
  OAI21_X1 U10405 ( .B1(n9377), .B2(n9332), .A(n9331), .ZN(n9333) );
  AOI21_X1 U10406 ( .B1(n9334), .B2(n9353), .A(n9333), .ZN(n9335) );
  OAI21_X1 U10407 ( .B1(n9336), .B2(n9355), .A(n9335), .ZN(P2_U3169) );
  INV_X1 U10408 ( .A(n9657), .ZN(n9771) );
  OAI211_X1 U10409 ( .C1(n9339), .C2(n9338), .A(n9337), .B(n5658), .ZN(n9344)
         );
  INV_X1 U10410 ( .A(n9340), .ZN(n9656) );
  AOI22_X1 U10411 ( .A1(n9380), .A2(n5193), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n9341) );
  OAI21_X1 U10412 ( .B1(n9655), .B2(n9376), .A(n9341), .ZN(n9342) );
  AOI21_X1 U10413 ( .B1(n9656), .B2(n9364), .A(n9342), .ZN(n9343) );
  OAI211_X1 U10414 ( .C1(n9771), .C2(n9383), .A(n9344), .B(n9343), .ZN(
        P2_U3173) );
  INV_X1 U10415 ( .A(n9345), .ZN(n9346) );
  AOI21_X1 U10416 ( .B1(n9348), .B2(n9347), .A(n9346), .ZN(n9356) );
  OAI22_X1 U10417 ( .A1(n9376), .A2(n9654), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9349), .ZN(n9350) );
  AOI21_X1 U10418 ( .B1(n9380), .B2(n9622), .A(n9350), .ZN(n9351) );
  OAI21_X1 U10419 ( .B1(n9624), .B2(n9377), .A(n9351), .ZN(n9352) );
  AOI21_X1 U10420 ( .B1(n9714), .B2(n9353), .A(n9352), .ZN(n9354) );
  OAI21_X1 U10421 ( .B1(n9356), .B2(n9355), .A(n9354), .ZN(P2_U3175) );
  OAI211_X1 U10422 ( .C1(n9359), .C2(n9358), .A(n9357), .B(n5658), .ZN(n9367)
         );
  INV_X1 U10423 ( .A(n9360), .ZN(n9365) );
  OAI22_X1 U10424 ( .A1(n9362), .A2(n9361), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9515), .ZN(n9363) );
  AOI21_X1 U10425 ( .B1(n9365), .B2(n9364), .A(n9363), .ZN(n9366) );
  OAI211_X1 U10426 ( .C1(n9780), .C2(n9383), .A(n9367), .B(n9366), .ZN(
        P2_U3178) );
  AOI22_X1 U10427 ( .A1(n9370), .A2(n9369), .B1(n9602), .B2(n9368), .ZN(n9374)
         );
  INV_X1 U10428 ( .A(n9371), .ZN(n9373) );
  OAI211_X1 U10429 ( .C1(n9374), .C2(n9373), .A(n5658), .B(n9372), .ZN(n9382)
         );
  OAI22_X1 U10430 ( .A1(n9376), .A2(n9602), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9375), .ZN(n9379) );
  NOR2_X1 U10431 ( .A1(n9377), .A2(n9577), .ZN(n9378) );
  AOI211_X1 U10432 ( .C1(n9380), .C2(n9385), .A(n9379), .B(n9378), .ZN(n9381)
         );
  OAI211_X1 U10433 ( .C1(n9756), .C2(n9383), .A(n9382), .B(n9381), .ZN(
        P2_U3180) );
  MUX2_X1 U10434 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n9535), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10435 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n9384), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10436 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9385), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10437 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n9386), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10438 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9387), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10439 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9612), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10440 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n9622), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U10441 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9611), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10442 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n5193), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10443 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9669), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10444 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9388), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10445 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9666), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10446 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9389), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10447 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9390), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10448 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9391), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10449 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n9392), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10450 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n9393), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10451 ( .A(n9394), .B(P2_DATAO_REG_12__SCAN_IN), .S(n10657), .Z(
        P2_U3503) );
  MUX2_X1 U10452 ( .A(n9395), .B(P2_DATAO_REG_11__SCAN_IN), .S(n10657), .Z(
        P2_U3502) );
  MUX2_X1 U10453 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n9396), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10454 ( .A(n9397), .B(P2_DATAO_REG_8__SCAN_IN), .S(n10657), .Z(
        P2_U3499) );
  MUX2_X1 U10455 ( .A(n9398), .B(P2_DATAO_REG_7__SCAN_IN), .S(n10657), .Z(
        P2_U3498) );
  MUX2_X1 U10456 ( .A(n9399), .B(P2_DATAO_REG_6__SCAN_IN), .S(n10657), .Z(
        P2_U3497) );
  MUX2_X1 U10457 ( .A(n9400), .B(P2_DATAO_REG_5__SCAN_IN), .S(n10657), .Z(
        P2_U3496) );
  MUX2_X1 U10458 ( .A(n9401), .B(P2_DATAO_REG_4__SCAN_IN), .S(n10657), .Z(
        P2_U3495) );
  MUX2_X1 U10459 ( .A(n9402), .B(P2_DATAO_REG_3__SCAN_IN), .S(n10657), .Z(
        P2_U3494) );
  MUX2_X1 U10460 ( .A(n9403), .B(P2_DATAO_REG_2__SCAN_IN), .S(n10657), .Z(
        P2_U3493) );
  MUX2_X1 U10461 ( .A(n9404), .B(P2_DATAO_REG_1__SCAN_IN), .S(n10657), .Z(
        P2_U3492) );
  MUX2_X1 U10462 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n9405), .S(P2_U3893), .Z(
        P2_U3491) );
  AOI21_X1 U10463 ( .B1(n9408), .B2(n9407), .A(n9406), .ZN(n9423) );
  INV_X1 U10464 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n9415) );
  OAI21_X1 U10465 ( .B1(n9411), .B2(n9410), .A(n9409), .ZN(n9412) );
  NAND2_X1 U10466 ( .A1(n9412), .A2(n10729), .ZN(n9414) );
  OAI211_X1 U10467 ( .C1(n10734), .C2(n9415), .A(n9414), .B(n9413), .ZN(n9420)
         );
  AOI21_X1 U10468 ( .B1(n5170), .B2(n9417), .A(n9416), .ZN(n9418) );
  NOR2_X1 U10469 ( .A1(n9418), .A2(n10717), .ZN(n9419) );
  AOI211_X1 U10470 ( .C1(n10722), .C2(n9421), .A(n9420), .B(n9419), .ZN(n9422)
         );
  OAI21_X1 U10471 ( .B1(n9423), .B2(n10724), .A(n9422), .ZN(P2_U3194) );
  INV_X1 U10472 ( .A(n10724), .ZN(n9517) );
  NOR2_X1 U10473 ( .A1(n9424), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9425) );
  OR2_X1 U10474 ( .A1(n9426), .A2(n9425), .ZN(n9428) );
  AOI21_X1 U10475 ( .B1(n9517), .B2(n9428), .A(n9427), .ZN(n9435) );
  NAND2_X1 U10476 ( .A1(n9505), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n9434) );
  OAI21_X1 U10477 ( .B1(n9431), .B2(n9430), .A(n9429), .ZN(n9432) );
  NAND2_X1 U10478 ( .A1(n9432), .A2(n10729), .ZN(n9433) );
  NAND3_X1 U10479 ( .A1(n9435), .A2(n9434), .A3(n9433), .ZN(n9441) );
  AOI21_X1 U10480 ( .B1(n9438), .B2(n9437), .A(n9436), .ZN(n9439) );
  NOR2_X1 U10481 ( .A1(n9439), .A2(n10717), .ZN(n9440) );
  AOI211_X1 U10482 ( .C1(n10722), .C2(n9442), .A(n9441), .B(n9440), .ZN(n9443)
         );
  INV_X1 U10483 ( .A(n9443), .ZN(P2_U3195) );
  AOI21_X1 U10484 ( .B1(n5173), .B2(n9445), .A(n9444), .ZN(n9459) );
  OAI21_X1 U10485 ( .B1(n9448), .B2(n9447), .A(n9446), .ZN(n9457) );
  NOR2_X1 U10486 ( .A1(n9521), .A2(n9449), .ZN(n9456) );
  AOI21_X1 U10487 ( .B1(n5122), .B2(n9451), .A(n9450), .ZN(n9454) );
  NAND2_X1 U10488 ( .A1(n9505), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n9453) );
  OAI211_X1 U10489 ( .C1(n9454), .C2(n10724), .A(n9453), .B(n9452), .ZN(n9455)
         );
  AOI211_X1 U10490 ( .C1(n10729), .C2(n9457), .A(n9456), .B(n9455), .ZN(n9458)
         );
  OAI21_X1 U10491 ( .B1(n9459), .B2(n10717), .A(n9458), .ZN(P2_U3196) );
  AOI21_X1 U10492 ( .B1(n9462), .B2(n9461), .A(n9460), .ZN(n9477) );
  OAI21_X1 U10493 ( .B1(n9465), .B2(n9464), .A(n9463), .ZN(n9475) );
  NOR2_X1 U10494 ( .A1(n9521), .A2(n9466), .ZN(n9474) );
  AOI21_X1 U10495 ( .B1(n9469), .B2(n9468), .A(n9467), .ZN(n9472) );
  NAND2_X1 U10496 ( .A1(n9505), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n9471) );
  OAI211_X1 U10497 ( .C1(n9472), .C2(n10724), .A(n9471), .B(n9470), .ZN(n9473)
         );
  AOI211_X1 U10498 ( .C1(n10729), .C2(n9475), .A(n9474), .B(n9473), .ZN(n9476)
         );
  OAI21_X1 U10499 ( .B1(n9477), .B2(n10717), .A(n9476), .ZN(P2_U3197) );
  AOI21_X1 U10500 ( .B1(n9480), .B2(n9479), .A(n9478), .ZN(n9495) );
  OAI21_X1 U10501 ( .B1(n9483), .B2(n9482), .A(n9481), .ZN(n9484) );
  NAND2_X1 U10502 ( .A1(n9484), .A2(n10729), .ZN(n9485) );
  OAI211_X1 U10503 ( .C1(n10734), .C2(n9487), .A(n9486), .B(n9485), .ZN(n9492)
         );
  AOI21_X1 U10504 ( .B1(n5165), .B2(n9489), .A(n9488), .ZN(n9490) );
  NOR2_X1 U10505 ( .A1(n9490), .A2(n10724), .ZN(n9491) );
  AOI211_X1 U10506 ( .C1(n10722), .C2(n9493), .A(n9492), .B(n9491), .ZN(n9494)
         );
  OAI21_X1 U10507 ( .B1(n9495), .B2(n10717), .A(n9494), .ZN(P2_U3198) );
  AOI21_X1 U10508 ( .B1(n9498), .B2(n9497), .A(n9496), .ZN(n9508) );
  XNOR2_X1 U10509 ( .A(n9500), .B(n9499), .ZN(n9507) );
  OAI21_X1 U10510 ( .B1(n10724), .B2(n9503), .A(n9502), .ZN(n9504) );
  AOI21_X1 U10511 ( .B1(n9510), .B2(n9509), .A(n5128), .ZN(n9532) );
  NOR2_X1 U10512 ( .A1(n9512), .A2(n9511), .ZN(n9514) );
  NOR2_X1 U10513 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9515), .ZN(n9516) );
  AOI21_X1 U10514 ( .B1(n9517), .B2(n5709), .A(n9516), .ZN(n9530) );
  INV_X1 U10515 ( .A(n9518), .ZN(n9520) );
  NAND2_X1 U10516 ( .A1(n9520), .A2(n9519), .ZN(n9523) );
  OAI21_X1 U10517 ( .B1(n9523), .B2(n10657), .A(n9521), .ZN(n9528) );
  NAND3_X1 U10518 ( .A1(n9523), .A2(n10729), .A3(n9522), .ZN(n9525) );
  INV_X1 U10519 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9524) );
  NAND2_X1 U10520 ( .A1(n9525), .A2(n5729), .ZN(n9526) );
  OAI21_X1 U10521 ( .B1(n9532), .B2(n10717), .A(n9531), .ZN(P2_U3200) );
  NOR2_X1 U10522 ( .A1(n9590), .A2(n9533), .ZN(n9540) );
  NOR2_X1 U10523 ( .A1(n9673), .A2(n9540), .ZN(n9536) );
  NAND2_X1 U10524 ( .A1(n9535), .A2(n9534), .ZN(n9739) );
  NAND2_X1 U10525 ( .A1(n9536), .A2(n9739), .ZN(n9538) );
  OAI21_X1 U10526 ( .B1(n10874), .B2(P2_REG2_REG_31__SCAN_IN), .A(n9538), .ZN(
        n9537) );
  OAI21_X1 U10527 ( .B1(n9741), .B2(n9647), .A(n9537), .ZN(P2_U3202) );
  OAI21_X1 U10528 ( .B1(n10874), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9538), .ZN(
        n9539) );
  OAI21_X1 U10529 ( .B1(n9744), .B2(n9647), .A(n9539), .ZN(P2_U3203) );
  AOI21_X1 U10530 ( .B1(n9673), .B2(P2_REG2_REG_29__SCAN_IN), .A(n9540), .ZN(
        n9541) );
  OAI21_X1 U10531 ( .B1(n9542), .B2(n9647), .A(n9541), .ZN(n9543) );
  AOI21_X1 U10532 ( .B1(n9545), .B2(n9544), .A(n9543), .ZN(n9546) );
  OAI21_X1 U10533 ( .B1(n9547), .B2(n9673), .A(n9546), .ZN(P2_U3204) );
  XNOR2_X1 U10534 ( .A(n9549), .B(n9548), .ZN(n9553) );
  AOI21_X1 U10535 ( .B1(n10871), .B2(n9554), .A(n9687), .ZN(n9560) );
  AOI22_X1 U10536 ( .A1(n9555), .A2(n10869), .B1(n9673), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n9559) );
  XNOR2_X1 U10537 ( .A(n9557), .B(n9556), .ZN(n9685) );
  NAND2_X1 U10538 ( .A1(n9685), .A2(n9677), .ZN(n9558) );
  OAI211_X1 U10539 ( .C1(n9560), .C2(n9673), .A(n9559), .B(n9558), .ZN(
        P2_U3205) );
  INV_X1 U10540 ( .A(n9690), .ZN(n9573) );
  XNOR2_X1 U10541 ( .A(n9567), .B(n9566), .ZN(n9691) );
  INV_X1 U10542 ( .A(n9568), .ZN(n9569) );
  AOI22_X1 U10543 ( .A1(n9673), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n10871), 
        .B2(n9569), .ZN(n9570) );
  OAI21_X1 U10544 ( .B1(n9752), .B2(n9647), .A(n9570), .ZN(n9571) );
  AOI21_X1 U10545 ( .B1(n9691), .B2(n9677), .A(n9571), .ZN(n9572) );
  OAI21_X1 U10546 ( .B1(n9573), .B2(n9673), .A(n9572), .ZN(P2_U3206) );
  XNOR2_X1 U10547 ( .A(n9574), .B(n9579), .ZN(n9575) );
  OAI222_X1 U10548 ( .A1(n9635), .A2(n9602), .B1(n9637), .B2(n9576), .C1(n9575), .C2(n9653), .ZN(n9695) );
  INV_X1 U10549 ( .A(n9695), .ZN(n9586) );
  INV_X1 U10550 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9578) );
  OAI22_X1 U10551 ( .A1(n10874), .A2(n9578), .B1(n9577), .B2(n9590), .ZN(n9583) );
  NOR2_X1 U10552 ( .A1(n9580), .A2(n9579), .ZN(n9694) );
  INV_X1 U10553 ( .A(n9696), .ZN(n9581) );
  NOR3_X1 U10554 ( .A1(n9694), .A2(n9581), .A3(n9629), .ZN(n9582) );
  AOI211_X1 U10555 ( .C1(n10869), .C2(n9584), .A(n9583), .B(n9582), .ZN(n9585)
         );
  OAI21_X1 U10556 ( .B1(n9586), .B2(n9673), .A(n9585), .ZN(P2_U3207) );
  XNOR2_X1 U10557 ( .A(n5149), .B(n9594), .ZN(n9587) );
  OAI222_X1 U10558 ( .A1(n9637), .A2(n9589), .B1(n9635), .B2(n9588), .C1(n9653), .C2(n9587), .ZN(n9701) );
  OAI22_X1 U10559 ( .A1(n9760), .A2(n9592), .B1(n9591), .B2(n9590), .ZN(n9593)
         );
  OAI21_X1 U10560 ( .B1(n9701), .B2(n9593), .A(n10874), .ZN(n9598) );
  NOR2_X1 U10561 ( .A1(n9595), .A2(n9594), .ZN(n9700) );
  NOR2_X1 U10562 ( .A1(n9700), .A2(n9629), .ZN(n9596) );
  AOI22_X1 U10563 ( .A1(n9596), .A2(n9702), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9673), .ZN(n9597) );
  NAND2_X1 U10564 ( .A1(n9598), .A2(n9597), .ZN(P2_U3208) );
  XOR2_X1 U10565 ( .A(n9604), .B(n9599), .Z(n9600) );
  OAI222_X1 U10566 ( .A1(n9637), .A2(n9602), .B1(n9635), .B2(n9601), .C1(n9600), .C2(n9653), .ZN(n9706) );
  INV_X1 U10567 ( .A(n9706), .ZN(n9609) );
  XOR2_X1 U10568 ( .A(n9604), .B(n9603), .Z(n9707) );
  AOI22_X1 U10569 ( .A1(n9673), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n10871), 
        .B2(n9605), .ZN(n9606) );
  OAI21_X1 U10570 ( .B1(n9764), .B2(n9647), .A(n9606), .ZN(n9607) );
  AOI21_X1 U10571 ( .B1(n9707), .B2(n9677), .A(n9607), .ZN(n9608) );
  OAI21_X1 U10572 ( .B1(n9609), .B2(n9673), .A(n9608), .ZN(P2_U3209) );
  XOR2_X1 U10573 ( .A(n9614), .B(n9610), .Z(n9613) );
  AOI222_X1 U10574 ( .A1(n9664), .A2(n9613), .B1(n9612), .B2(n9668), .C1(n9611), .C2(n9667), .ZN(n9713) );
  XOR2_X1 U10575 ( .A(n9615), .B(n9614), .Z(n9711) );
  AOI22_X1 U10576 ( .A1(n9673), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n10871), 
        .B2(n9616), .ZN(n9617) );
  OAI21_X1 U10577 ( .B1(n9618), .B2(n9647), .A(n9617), .ZN(n9619) );
  AOI21_X1 U10578 ( .B1(n9711), .B2(n9677), .A(n9619), .ZN(n9620) );
  OAI21_X1 U10579 ( .B1(n9713), .B2(n9673), .A(n9620), .ZN(P2_U3210) );
  XNOR2_X1 U10580 ( .A(n9621), .B(n9627), .ZN(n9623) );
  AOI222_X1 U10581 ( .A1(n9664), .A2(n9623), .B1(n9622), .B2(n9668), .C1(n5193), .C2(n9667), .ZN(n9716) );
  INV_X1 U10582 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n9625) );
  OAI22_X1 U10583 ( .A1(n10874), .A2(n9625), .B1(n9624), .B2(n9590), .ZN(n9631) );
  OAI21_X1 U10584 ( .B1(n9628), .B2(n9627), .A(n9626), .ZN(n9717) );
  NOR2_X1 U10585 ( .A1(n9717), .A2(n9629), .ZN(n9630) );
  AOI211_X1 U10586 ( .C1(n10869), .C2(n9714), .A(n9631), .B(n9630), .ZN(n9632)
         );
  OAI21_X1 U10587 ( .B1(n9716), .B2(n9673), .A(n9632), .ZN(P2_U3211) );
  XNOR2_X1 U10588 ( .A(n9633), .B(n9634), .ZN(n9640) );
  OAI22_X1 U10589 ( .A1(n9638), .A2(n9637), .B1(n9636), .B2(n9635), .ZN(n9639)
         );
  AOI21_X1 U10590 ( .B1(n9640), .B2(n9664), .A(n9639), .ZN(n9723) );
  OR2_X1 U10591 ( .A1(n9642), .A2(n9641), .ZN(n9643) );
  AND2_X1 U10592 ( .A1(n9644), .A2(n9643), .ZN(n9721) );
  AOI22_X1 U10593 ( .A1(n9673), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n10871), 
        .B2(n9645), .ZN(n9646) );
  OAI21_X1 U10594 ( .B1(n9648), .B2(n9647), .A(n9646), .ZN(n9649) );
  AOI21_X1 U10595 ( .B1(n9721), .B2(n9677), .A(n9649), .ZN(n9650) );
  OAI21_X1 U10596 ( .B1(n9723), .B2(n9673), .A(n9650), .ZN(P2_U3212) );
  AOI21_X1 U10597 ( .B1(n9659), .B2(n9651), .A(n5174), .ZN(n9652) );
  OAI222_X1 U10598 ( .A1(n9635), .A2(n9655), .B1(n9637), .B2(n9654), .C1(n9653), .C2(n9652), .ZN(n9724) );
  AOI21_X1 U10599 ( .B1(n10871), .B2(n9656), .A(n9724), .ZN(n9662) );
  AOI22_X1 U10600 ( .A1(n9657), .A2(n10869), .B1(P2_REG2_REG_20__SCAN_IN), 
        .B2(n9673), .ZN(n9661) );
  XNOR2_X1 U10601 ( .A(n9658), .B(n9659), .ZN(n9725) );
  NAND2_X1 U10602 ( .A1(n9725), .A2(n9677), .ZN(n9660) );
  OAI211_X1 U10603 ( .C1(n9662), .C2(n9673), .A(n9661), .B(n9660), .ZN(
        P2_U3213) );
  OAI211_X1 U10604 ( .C1(n9665), .C2(n6330), .A(n9664), .B(n9663), .ZN(n9671)
         );
  AOI22_X1 U10605 ( .A1(n9669), .A2(n9668), .B1(n9667), .B2(n9666), .ZN(n9670)
         );
  NAND2_X1 U10606 ( .A1(n9671), .A2(n9670), .ZN(n9728) );
  AOI21_X1 U10607 ( .B1(n10871), .B2(n9672), .A(n9728), .ZN(n9680) );
  AOI22_X1 U10608 ( .A1(n9674), .A2(n10869), .B1(P2_REG2_REG_19__SCAN_IN), 
        .B2(n9673), .ZN(n9679) );
  XNOR2_X1 U10609 ( .A(n9675), .B(n9676), .ZN(n9729) );
  NAND2_X1 U10610 ( .A1(n9729), .A2(n9677), .ZN(n9678) );
  OAI211_X1 U10611 ( .C1(n9680), .C2(n9673), .A(n9679), .B(n9678), .ZN(
        P2_U3214) );
  NOR2_X1 U10612 ( .A1(n9683), .A2(n9739), .ZN(n9682) );
  AOI21_X1 U10613 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n9683), .A(n9682), .ZN(
        n9681) );
  OAI21_X1 U10614 ( .B1(n9741), .B2(n9738), .A(n9681), .ZN(P2_U3490) );
  AOI21_X1 U10615 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n9683), .A(n9682), .ZN(
        n9684) );
  OAI21_X1 U10616 ( .B1(n9744), .B2(n9738), .A(n9684), .ZN(P2_U3489) );
  MUX2_X1 U10617 ( .A(n9688), .B(n9745), .S(n9735), .Z(n9689) );
  OAI21_X1 U10618 ( .B1(n9748), .B2(n9738), .A(n9689), .ZN(P2_U3487) );
  AOI21_X1 U10619 ( .B1(n9733), .B2(n9691), .A(n9690), .ZN(n9749) );
  MUX2_X1 U10620 ( .A(n9692), .B(n9749), .S(n9735), .Z(n9693) );
  OAI21_X1 U10621 ( .B1(n9752), .B2(n9738), .A(n9693), .ZN(P2_U3486) );
  NOR2_X1 U10622 ( .A1(n9694), .A2(n9718), .ZN(n9697) );
  AOI21_X1 U10623 ( .B1(n9697), .B2(n9696), .A(n9695), .ZN(n9753) );
  MUX2_X1 U10624 ( .A(n9698), .B(n9753), .S(n9735), .Z(n9699) );
  OAI21_X1 U10625 ( .B1(n9756), .B2(n9738), .A(n9699), .ZN(P2_U3485) );
  NOR2_X1 U10626 ( .A1(n9700), .A2(n9718), .ZN(n9703) );
  AOI21_X1 U10627 ( .B1(n9703), .B2(n9702), .A(n9701), .ZN(n9757) );
  MUX2_X1 U10628 ( .A(n9704), .B(n9757), .S(n9735), .Z(n9705) );
  OAI21_X1 U10629 ( .B1(n9760), .B2(n9738), .A(n9705), .ZN(P2_U3484) );
  AOI21_X1 U10630 ( .B1(n9733), .B2(n9707), .A(n9706), .ZN(n9761) );
  MUX2_X1 U10631 ( .A(n9708), .B(n9761), .S(n9735), .Z(n9709) );
  OAI21_X1 U10632 ( .B1(n9764), .B2(n9738), .A(n9709), .ZN(P2_U3483) );
  AOI22_X1 U10633 ( .A1(n9711), .A2(n9733), .B1(n9720), .B2(n9710), .ZN(n9712)
         );
  NAND2_X1 U10634 ( .A1(n9713), .A2(n9712), .ZN(n9765) );
  MUX2_X1 U10635 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9765), .S(n9735), .Z(
        P2_U3482) );
  NAND2_X1 U10636 ( .A1(n9714), .A2(n9720), .ZN(n9715) );
  OAI211_X1 U10637 ( .C1(n9718), .C2(n9717), .A(n9716), .B(n9715), .ZN(n9766)
         );
  MUX2_X1 U10638 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9766), .S(n9735), .Z(
        P2_U3481) );
  AOI22_X1 U10639 ( .A1(n9721), .A2(n9733), .B1(n9720), .B2(n9719), .ZN(n9722)
         );
  NAND2_X1 U10640 ( .A1(n9723), .A2(n9722), .ZN(n9767) );
  MUX2_X1 U10641 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9767), .S(n9735), .Z(
        P2_U3480) );
  AOI21_X1 U10642 ( .B1(n9725), .B2(n9733), .A(n9724), .ZN(n9768) );
  MUX2_X1 U10643 ( .A(n9726), .B(n9768), .S(n9735), .Z(n9727) );
  OAI21_X1 U10644 ( .B1(n9771), .B2(n9738), .A(n9727), .ZN(P2_U3479) );
  AOI21_X1 U10645 ( .B1(n9729), .B2(n9733), .A(n9728), .ZN(n9772) );
  MUX2_X1 U10646 ( .A(n9730), .B(n9772), .S(n9735), .Z(n9731) );
  OAI21_X1 U10647 ( .B1(n9775), .B2(n9738), .A(n9731), .ZN(P2_U3478) );
  AOI21_X1 U10648 ( .B1(n9734), .B2(n9733), .A(n9732), .ZN(n9776) );
  MUX2_X1 U10649 ( .A(n9736), .B(n9776), .S(n9735), .Z(n9737) );
  OAI21_X1 U10650 ( .B1(n9780), .B2(n9738), .A(n9737), .ZN(P2_U3477) );
  NOR2_X1 U10651 ( .A1(n11015), .A2(n9739), .ZN(n9742) );
  AOI21_X1 U10652 ( .B1(P2_REG0_REG_31__SCAN_IN), .B2(n11015), .A(n9742), .ZN(
        n9740) );
  OAI21_X1 U10653 ( .B1(n9741), .B2(n9779), .A(n9740), .ZN(P2_U3458) );
  AOI21_X1 U10654 ( .B1(P2_REG0_REG_30__SCAN_IN), .B2(n11015), .A(n9742), .ZN(
        n9743) );
  OAI21_X1 U10655 ( .B1(n9744), .B2(n9779), .A(n9743), .ZN(P2_U3457) );
  MUX2_X1 U10656 ( .A(n9746), .B(n9745), .S(n11017), .Z(n9747) );
  OAI21_X1 U10657 ( .B1(n9748), .B2(n9779), .A(n9747), .ZN(P2_U3455) );
  MUX2_X1 U10658 ( .A(n9750), .B(n9749), .S(n11017), .Z(n9751) );
  OAI21_X1 U10659 ( .B1(n9752), .B2(n9779), .A(n9751), .ZN(P2_U3454) );
  MUX2_X1 U10660 ( .A(n9754), .B(n9753), .S(n11017), .Z(n9755) );
  OAI21_X1 U10661 ( .B1(n9756), .B2(n9779), .A(n9755), .ZN(P2_U3453) );
  MUX2_X1 U10662 ( .A(n9758), .B(n9757), .S(n11017), .Z(n9759) );
  OAI21_X1 U10663 ( .B1(n9760), .B2(n9779), .A(n9759), .ZN(P2_U3452) );
  MUX2_X1 U10664 ( .A(n9762), .B(n9761), .S(n11017), .Z(n9763) );
  OAI21_X1 U10665 ( .B1(n9764), .B2(n9779), .A(n9763), .ZN(P2_U3451) );
  MUX2_X1 U10666 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9765), .S(n11017), .Z(
        P2_U3450) );
  MUX2_X1 U10667 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9766), .S(n11017), .Z(
        P2_U3449) );
  MUX2_X1 U10668 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9767), .S(n11017), .Z(
        P2_U3448) );
  MUX2_X1 U10669 ( .A(n9769), .B(n9768), .S(n11017), .Z(n9770) );
  OAI21_X1 U10670 ( .B1(n9771), .B2(n9779), .A(n9770), .ZN(P2_U3447) );
  MUX2_X1 U10671 ( .A(n9773), .B(n9772), .S(n11017), .Z(n9774) );
  OAI21_X1 U10672 ( .B1(n9775), .B2(n9779), .A(n9774), .ZN(P2_U3446) );
  MUX2_X1 U10673 ( .A(n9777), .B(n9776), .S(n11017), .Z(n9778) );
  OAI21_X1 U10674 ( .B1(n9780), .B2(n9779), .A(n9778), .ZN(P2_U3444) );
  INV_X1 U10675 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9782) );
  NAND3_X1 U10676 ( .A1(n9782), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n9785) );
  OAI22_X1 U10677 ( .A1(n9781), .A2(n9785), .B1(n9784), .B2(n9783), .ZN(n9786)
         );
  AOI21_X1 U10678 ( .B1(n7309), .B2(n9787), .A(n9786), .ZN(n9788) );
  INV_X1 U10679 ( .A(n9788), .ZN(P2_U3264) );
  AOI21_X1 U10680 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n9790), .A(n9789), .ZN(
        n9791) );
  OAI21_X1 U10681 ( .B1(n9793), .B2(n9792), .A(n9791), .ZN(P2_U3267) );
  MUX2_X1 U10682 ( .A(n9794), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10683 ( .A1(n9799), .A2(n9948), .ZN(n9796) );
  OR2_X1 U10684 ( .A1(n9924), .A2(n7808), .ZN(n9795) );
  NAND2_X1 U10685 ( .A1(n9796), .A2(n9795), .ZN(n9797) );
  XNOR2_X1 U10686 ( .A(n9797), .B(n9951), .ZN(n9804) );
  NOR2_X1 U10687 ( .A1(n9924), .A2(n9901), .ZN(n9798) );
  AOI21_X1 U10688 ( .B1(n9799), .B2(n9863), .A(n9798), .ZN(n9805) );
  XNOR2_X1 U10689 ( .A(n9804), .B(n9805), .ZN(n10037) );
  NAND2_X1 U10690 ( .A1(n9801), .A2(n9800), .ZN(n10035) );
  AND2_X1 U10691 ( .A1(n10037), .A2(n10035), .ZN(n9802) );
  INV_X1 U10692 ( .A(n9804), .ZN(n9806) );
  NAND2_X1 U10693 ( .A1(n10255), .A2(n9948), .ZN(n9808) );
  NAND2_X1 U10694 ( .A1(n10551), .A2(n9954), .ZN(n9807) );
  NAND2_X1 U10695 ( .A1(n9808), .A2(n9807), .ZN(n9809) );
  XNOR2_X1 U10696 ( .A(n9809), .B(n9951), .ZN(n9810) );
  AOI22_X1 U10697 ( .A1(n10255), .A2(n9954), .B1(n9953), .B2(n10551), .ZN(
        n9920) );
  INV_X1 U10698 ( .A(n9813), .ZN(n9814) );
  NAND2_X1 U10699 ( .A1(n10556), .A2(n9948), .ZN(n9816) );
  OR2_X1 U10700 ( .A1(n10465), .A2(n7808), .ZN(n9815) );
  NAND2_X1 U10701 ( .A1(n9816), .A2(n9815), .ZN(n9817) );
  XNOR2_X1 U10702 ( .A(n9817), .B(n9899), .ZN(n9823) );
  NOR2_X1 U10703 ( .A1(n10465), .A2(n9901), .ZN(n9818) );
  AOI21_X1 U10704 ( .B1(n10556), .B2(n9954), .A(n9818), .ZN(n10080) );
  NAND2_X1 U10705 ( .A1(n10480), .A2(n9948), .ZN(n9820) );
  OR2_X1 U10706 ( .A1(n10450), .A2(n7808), .ZN(n9819) );
  NAND2_X1 U10707 ( .A1(n9820), .A2(n9819), .ZN(n9821) );
  XNOR2_X1 U10708 ( .A(n9821), .B(n9899), .ZN(n9825) );
  NOR2_X1 U10709 ( .A1(n10450), .A2(n9901), .ZN(n9822) );
  AOI21_X1 U10710 ( .B1(n10480), .B2(n9954), .A(n9822), .ZN(n9824) );
  XNOR2_X1 U10711 ( .A(n9825), .B(n9824), .ZN(n9996) );
  INV_X1 U10712 ( .A(n10080), .ZN(n9997) );
  NOR2_X1 U10713 ( .A1(n10463), .A2(n7808), .ZN(n9826) );
  AOI21_X1 U10714 ( .B1(n10543), .B2(n9948), .A(n9826), .ZN(n9827) );
  XNOR2_X1 U10715 ( .A(n9827), .B(n9951), .ZN(n9831) );
  NOR2_X1 U10716 ( .A1(n10463), .A2(n9901), .ZN(n9828) );
  AOI21_X1 U10717 ( .B1(n10543), .B2(n9954), .A(n9828), .ZN(n9830) );
  NOR2_X1 U10718 ( .A1(n9831), .A2(n9830), .ZN(n10008) );
  NAND2_X1 U10719 ( .A1(n10005), .A2(n9829), .ZN(n9832) );
  NAND2_X1 U10720 ( .A1(n9831), .A2(n9830), .ZN(n10006) );
  NAND2_X1 U10721 ( .A1(n9832), .A2(n10006), .ZN(n9937) );
  NAND2_X1 U10722 ( .A1(n10428), .A2(n9948), .ZN(n9834) );
  OR2_X1 U10723 ( .A1(n10433), .A2(n7808), .ZN(n9833) );
  NAND2_X1 U10724 ( .A1(n9834), .A2(n9833), .ZN(n9835) );
  XNOR2_X1 U10725 ( .A(n9835), .B(n9951), .ZN(n9940) );
  NOR2_X1 U10726 ( .A1(n10433), .A2(n9901), .ZN(n9836) );
  AOI21_X1 U10727 ( .B1(n10428), .B2(n9954), .A(n9836), .ZN(n9939) );
  INV_X1 U10728 ( .A(n9939), .ZN(n9842) );
  NAND2_X1 U10729 ( .A1(n10260), .A2(n9954), .ZN(n9838) );
  NAND2_X1 U10730 ( .A1(n10417), .A2(n9953), .ZN(n9837) );
  NAND2_X1 U10731 ( .A1(n10260), .A2(n9948), .ZN(n9840) );
  NAND2_X1 U10732 ( .A1(n10417), .A2(n9954), .ZN(n9839) );
  NAND2_X1 U10733 ( .A1(n9840), .A2(n9839), .ZN(n9841) );
  XNOR2_X1 U10734 ( .A(n9841), .B(n9899), .ZN(n9938) );
  INV_X1 U10735 ( .A(n9938), .ZN(n9845) );
  AOI22_X1 U10736 ( .A1(n9940), .A2(n9842), .B1(n10058), .B2(n9845), .ZN(n9848) );
  AOI21_X1 U10737 ( .B1(n9938), .B2(n9843), .A(n9939), .ZN(n9846) );
  NAND2_X1 U10738 ( .A1(n9939), .A2(n9843), .ZN(n9844) );
  OAI22_X1 U10739 ( .A1(n9846), .A2(n9940), .B1(n9845), .B2(n9844), .ZN(n9847)
         );
  NAND2_X1 U10740 ( .A1(n10537), .A2(n9948), .ZN(n9850) );
  OR2_X1 U10741 ( .A1(n10262), .A2(n7808), .ZN(n9849) );
  NAND2_X1 U10742 ( .A1(n9850), .A2(n9849), .ZN(n9851) );
  XNOR2_X1 U10743 ( .A(n9851), .B(n9951), .ZN(n9853) );
  OAI22_X1 U10744 ( .A1(n10407), .A2(n7808), .B1(n10262), .B2(n9901), .ZN(
        n9852) );
  XNOR2_X1 U10745 ( .A(n9853), .B(n9852), .ZN(n10026) );
  NAND2_X1 U10746 ( .A1(n10531), .A2(n9948), .ZN(n9855) );
  OR2_X1 U10747 ( .A1(n10263), .A2(n7808), .ZN(n9854) );
  NAND2_X1 U10748 ( .A1(n9855), .A2(n9854), .ZN(n9856) );
  XNOR2_X1 U10749 ( .A(n9856), .B(n9899), .ZN(n9859) );
  NOR2_X1 U10750 ( .A1(n10263), .A2(n9901), .ZN(n9857) );
  AOI21_X1 U10751 ( .B1(n10531), .B2(n9954), .A(n9857), .ZN(n9858) );
  OR2_X1 U10752 ( .A1(n9859), .A2(n9858), .ZN(n9973) );
  NAND2_X1 U10753 ( .A1(n9859), .A2(n9858), .ZN(n9972) );
  OAI22_X1 U10754 ( .A1(n10376), .A2(n9860), .B1(n10264), .B2(n7808), .ZN(
        n9861) );
  XOR2_X1 U10755 ( .A(n9951), .B(n9861), .Z(n9864) );
  NOR2_X1 U10756 ( .A1(n10264), .A2(n9901), .ZN(n9862) );
  AOI21_X1 U10757 ( .B1(n10525), .B2(n9863), .A(n9862), .ZN(n10049) );
  NAND2_X1 U10758 ( .A1(n9865), .A2(n9864), .ZN(n10047) );
  NAND2_X1 U10759 ( .A1(n10520), .A2(n9948), .ZN(n9867) );
  NAND2_X1 U10760 ( .A1(n10380), .A2(n9954), .ZN(n9866) );
  NAND2_X1 U10761 ( .A1(n9867), .A2(n9866), .ZN(n9868) );
  XNOR2_X1 U10762 ( .A(n9868), .B(n9951), .ZN(n9872) );
  NAND2_X1 U10763 ( .A1(n10520), .A2(n9954), .ZN(n9870) );
  NAND2_X1 U10764 ( .A1(n10380), .A2(n9953), .ZN(n9869) );
  NAND2_X1 U10765 ( .A1(n9870), .A2(n9869), .ZN(n9871) );
  AOI21_X1 U10766 ( .B1(n9872), .B2(n9871), .A(n10016), .ZN(n9931) );
  NAND2_X1 U10767 ( .A1(n9930), .A2(n9931), .ZN(n9929) );
  INV_X1 U10768 ( .A(n10016), .ZN(n9873) );
  NAND2_X1 U10769 ( .A1(n9929), .A2(n9873), .ZN(n9881) );
  NAND2_X1 U10770 ( .A1(n10514), .A2(n9948), .ZN(n9875) );
  OR2_X1 U10771 ( .A1(n9986), .A2(n7808), .ZN(n9874) );
  NAND2_X1 U10772 ( .A1(n9875), .A2(n9874), .ZN(n9876) );
  XNOR2_X1 U10773 ( .A(n9876), .B(n9899), .ZN(n9879) );
  NOR2_X1 U10774 ( .A1(n9986), .A2(n9901), .ZN(n9877) );
  AOI21_X1 U10775 ( .B1(n10514), .B2(n9954), .A(n9877), .ZN(n9878) );
  NAND2_X1 U10776 ( .A1(n9879), .A2(n9878), .ZN(n9882) );
  OR2_X1 U10777 ( .A1(n9879), .A2(n9878), .ZN(n9880) );
  NAND2_X1 U10778 ( .A1(n9881), .A2(n10015), .ZN(n10018) );
  NAND2_X1 U10779 ( .A1(n10018), .A2(n9882), .ZN(n9983) );
  OAI22_X1 U10780 ( .A1(n5390), .A2(n7808), .B1(n10318), .B2(n9901), .ZN(n9890) );
  NAND2_X1 U10781 ( .A1(n10510), .A2(n9948), .ZN(n9884) );
  NAND2_X1 U10782 ( .A1(n10351), .A2(n9954), .ZN(n9883) );
  NAND2_X1 U10783 ( .A1(n9884), .A2(n9883), .ZN(n9885) );
  XNOR2_X1 U10784 ( .A(n9885), .B(n9951), .ZN(n9891) );
  XOR2_X1 U10785 ( .A(n9890), .B(n9891), .Z(n9984) );
  NAND2_X1 U10786 ( .A1(n10506), .A2(n9948), .ZN(n9887) );
  OR2_X1 U10787 ( .A1(n10305), .A2(n7808), .ZN(n9886) );
  NAND2_X1 U10788 ( .A1(n9887), .A2(n9886), .ZN(n9888) );
  XNOR2_X1 U10789 ( .A(n9888), .B(n9899), .ZN(n9893) );
  NOR2_X1 U10790 ( .A1(n10305), .A2(n9901), .ZN(n9889) );
  AOI21_X1 U10791 ( .B1(n10506), .B2(n9954), .A(n9889), .ZN(n9894) );
  XNOR2_X1 U10792 ( .A(n9893), .B(n9894), .ZN(n10066) );
  NOR2_X1 U10793 ( .A1(n9891), .A2(n9890), .ZN(n10067) );
  NOR2_X1 U10794 ( .A1(n10066), .A2(n10067), .ZN(n9892) );
  INV_X1 U10795 ( .A(n9893), .ZN(n9896) );
  INV_X1 U10796 ( .A(n9894), .ZN(n9895) );
  NAND2_X1 U10797 ( .A1(n9896), .A2(n9895), .ZN(n9908) );
  NAND2_X1 U10798 ( .A1(n10501), .A2(n9948), .ZN(n9898) );
  OR2_X1 U10799 ( .A1(n10319), .A2(n7808), .ZN(n9897) );
  NAND2_X1 U10800 ( .A1(n9898), .A2(n9897), .ZN(n9900) );
  XNOR2_X1 U10801 ( .A(n9900), .B(n9899), .ZN(n9904) );
  INV_X1 U10802 ( .A(n9904), .ZN(n9906) );
  NOR2_X1 U10803 ( .A1(n10319), .A2(n9901), .ZN(n9902) );
  AOI21_X1 U10804 ( .B1(n10501), .B2(n9954), .A(n9902), .ZN(n9903) );
  INV_X1 U10805 ( .A(n9903), .ZN(n9905) );
  AOI21_X1 U10806 ( .B1(n9906), .B2(n9905), .A(n9966), .ZN(n9907) );
  AOI21_X1 U10807 ( .B1(n10069), .B2(n9908), .A(n9907), .ZN(n9912) );
  INV_X1 U10808 ( .A(n9907), .ZN(n9910) );
  INV_X1 U10809 ( .A(n9908), .ZN(n9909) );
  NOR2_X1 U10810 ( .A1(n9910), .A2(n9909), .ZN(n9911) );
  AOI22_X1 U10811 ( .A1(n10087), .A2(n10271), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9916) );
  NOR2_X1 U10812 ( .A1(n10041), .A2(n10464), .ZN(n10072) );
  AOI22_X1 U10813 ( .A1(n10072), .A2(n9913), .B1(n10071), .B2(n10308), .ZN(
        n9915) );
  NAND2_X1 U10814 ( .A1(n10501), .A2(n10073), .ZN(n9914) );
  NAND4_X1 U10815 ( .A1(n9917), .A2(n9916), .A3(n9915), .A4(n9914), .ZN(
        P1_U3214) );
  OAI21_X1 U10816 ( .B1(n9920), .B2(n9919), .A(n9918), .ZN(n9921) );
  NAND2_X1 U10817 ( .A1(n9921), .A2(n10081), .ZN(n9928) );
  NAND2_X1 U10818 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n10119)
         );
  INV_X1 U10819 ( .A(n10119), .ZN(n9926) );
  INV_X1 U10820 ( .A(n10072), .ZN(n10085) );
  INV_X1 U10821 ( .A(n9922), .ZN(n9923) );
  OAI22_X1 U10822 ( .A1(n10085), .A2(n9924), .B1(n10084), .B2(n9923), .ZN(
        n9925) );
  AOI211_X1 U10823 ( .C1(n10087), .C2(n5693), .A(n9926), .B(n9925), .ZN(n9927)
         );
  OAI211_X1 U10824 ( .C1(n10975), .C2(n10090), .A(n9928), .B(n9927), .ZN(
        P1_U3215) );
  OAI21_X1 U10825 ( .B1(n9931), .B2(n9930), .A(n9929), .ZN(n9932) );
  NAND2_X1 U10826 ( .A1(n9932), .A2(n10081), .ZN(n9936) );
  INV_X1 U10827 ( .A(n9986), .ZN(n10363) );
  AOI22_X1 U10828 ( .A1(n10087), .A2(n10363), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9935) );
  INV_X1 U10829 ( .A(n10264), .ZN(n10389) );
  AOI22_X1 U10830 ( .A1(n10072), .A2(n10389), .B1(n10071), .B2(n10358), .ZN(
        n9934) );
  NAND2_X1 U10831 ( .A1(n10520), .A2(n10073), .ZN(n9933) );
  NAND4_X1 U10832 ( .A1(n9936), .A2(n9935), .A3(n9934), .A4(n9933), .ZN(
        P1_U3216) );
  XNOR2_X1 U10833 ( .A(n9937), .B(n9938), .ZN(n10059) );
  NOR2_X1 U10834 ( .A1(n10059), .A2(n10058), .ZN(n10057) );
  AOI21_X1 U10835 ( .B1(n9938), .B2(n9937), .A(n10057), .ZN(n9942) );
  XNOR2_X1 U10836 ( .A(n9940), .B(n9939), .ZN(n9941) );
  XNOR2_X1 U10837 ( .A(n9942), .B(n9941), .ZN(n9947) );
  AOI22_X1 U10838 ( .A1(n10072), .A2(n10417), .B1(n10071), .B2(n9943), .ZN(
        n9944) );
  NAND2_X1 U10839 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n10218)
         );
  OAI211_X1 U10840 ( .C1(n10061), .C2(n10262), .A(n9944), .B(n10218), .ZN(
        n9945) );
  AOI21_X1 U10841 ( .B1(n10428), .B2(n10073), .A(n9945), .ZN(n9946) );
  OAI21_X1 U10842 ( .B1(n9947), .B2(n10064), .A(n9946), .ZN(P1_U3219) );
  NAND2_X1 U10843 ( .A1(n10495), .A2(n9948), .ZN(n9950) );
  NAND2_X1 U10844 ( .A1(n10271), .A2(n9954), .ZN(n9949) );
  NAND2_X1 U10845 ( .A1(n9950), .A2(n9949), .ZN(n9952) );
  XNOR2_X1 U10846 ( .A(n9952), .B(n9951), .ZN(n9956) );
  AOI22_X1 U10847 ( .A1(n10495), .A2(n9954), .B1(n9953), .B2(n10271), .ZN(
        n9955) );
  XNOR2_X1 U10848 ( .A(n9956), .B(n9955), .ZN(n9967) );
  INV_X1 U10849 ( .A(n9967), .ZN(n9957) );
  NAND3_X1 U10850 ( .A1(n9958), .A2(n9957), .A3(n5730), .ZN(n9971) );
  NAND3_X1 U10851 ( .A1(n9959), .A2(n10081), .A3(n9967), .ZN(n9970) );
  INV_X1 U10852 ( .A(n10288), .ZN(n9964) );
  OR2_X1 U10853 ( .A1(n9960), .A2(n10462), .ZN(n9962) );
  OR2_X1 U10854 ( .A1(n10319), .A2(n10464), .ZN(n9961) );
  NAND2_X1 U10855 ( .A1(n9962), .A2(n9961), .ZN(n10293) );
  AOI22_X1 U10856 ( .A1(n10293), .A2(n10029), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9963) );
  OAI21_X1 U10857 ( .B1(n9964), .B2(n10084), .A(n9963), .ZN(n9965) );
  AOI21_X1 U10858 ( .B1(n10495), .B2(n10073), .A(n9965), .ZN(n9969) );
  NAND3_X1 U10859 ( .A1(n9967), .A2(n9966), .A3(n10081), .ZN(n9968) );
  NAND4_X1 U10860 ( .A1(n9971), .A2(n9970), .A3(n9969), .A4(n9968), .ZN(
        P1_U3220) );
  NAND2_X1 U10861 ( .A1(n9973), .A2(n9972), .ZN(n9974) );
  XNOR2_X1 U10862 ( .A(n9975), .B(n9974), .ZN(n9981) );
  INV_X1 U10863 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9976) );
  OAI22_X1 U10864 ( .A1(n10061), .A2(n10264), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9976), .ZN(n9979) );
  INV_X1 U10865 ( .A(n10394), .ZN(n9977) );
  OAI22_X1 U10866 ( .A1(n10085), .A2(n10262), .B1(n10084), .B2(n9977), .ZN(
        n9978) );
  AOI211_X1 U10867 ( .C1(n10531), .C2(n10073), .A(n9979), .B(n9978), .ZN(n9980) );
  OAI21_X1 U10868 ( .B1(n9981), .B2(n10064), .A(n9980), .ZN(P1_U3223) );
  OAI21_X1 U10869 ( .B1(n9984), .B2(n9983), .A(n9982), .ZN(n9985) );
  NAND2_X1 U10870 ( .A1(n9985), .A2(n10081), .ZN(n9992) );
  OR2_X1 U10871 ( .A1(n9986), .A2(n10464), .ZN(n9988) );
  OR2_X1 U10872 ( .A1(n10305), .A2(n10462), .ZN(n9987) );
  NAND2_X1 U10873 ( .A1(n9988), .A2(n9987), .ZN(n10336) );
  AOI22_X1 U10874 ( .A1(n10336), .A2(n10029), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9991) );
  NAND2_X1 U10875 ( .A1(n10510), .A2(n10073), .ZN(n9990) );
  NAND2_X1 U10876 ( .A1(n10071), .A2(n10331), .ZN(n9989) );
  NAND4_X1 U10877 ( .A1(n9992), .A2(n9991), .A3(n9990), .A4(n9989), .ZN(
        P1_U3225) );
  NOR2_X1 U10878 ( .A1(n5110), .A2(n9998), .ZN(n9993) );
  AOI21_X1 U10879 ( .B1(n5110), .B2(n9998), .A(n9993), .ZN(n10079) );
  NAND2_X1 U10880 ( .A1(n10079), .A2(n10080), .ZN(n10078) );
  INV_X1 U10881 ( .A(n9993), .ZN(n9994) );
  AND3_X1 U10882 ( .A1(n10078), .A2(n9996), .A3(n9994), .ZN(n10000) );
  AOI211_X1 U10883 ( .C1(n9998), .C2(n9997), .A(n9996), .B(n9995), .ZN(n9999)
         );
  OAI21_X1 U10884 ( .B1(n10000), .B2(n9999), .A(n10081), .ZN(n10004) );
  INV_X1 U10885 ( .A(n10463), .ZN(n10258) );
  AND2_X1 U10886 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10167) );
  INV_X1 U10887 ( .A(n10001), .ZN(n10473) );
  OAI22_X1 U10888 ( .A1(n10085), .A2(n10465), .B1(n10084), .B2(n10473), .ZN(
        n10002) );
  AOI211_X1 U10889 ( .C1(n10087), .C2(n10258), .A(n10167), .B(n10002), .ZN(
        n10003) );
  OAI211_X1 U10890 ( .C1(n11008), .C2(n10090), .A(n10004), .B(n10003), .ZN(
        P1_U3226) );
  INV_X1 U10891 ( .A(n10006), .ZN(n10007) );
  NOR2_X1 U10892 ( .A1(n10008), .A2(n10007), .ZN(n10009) );
  XNOR2_X1 U10893 ( .A(n10010), .B(n10009), .ZN(n10014) );
  INV_X1 U10894 ( .A(n10450), .ZN(n10553) );
  AOI22_X1 U10895 ( .A1(n10072), .A2(n10553), .B1(n10071), .B2(n10453), .ZN(
        n10011) );
  NAND2_X1 U10896 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10185)
         );
  OAI211_X1 U10897 ( .C1(n10061), .C2(n10451), .A(n10011), .B(n10185), .ZN(
        n10012) );
  AOI21_X1 U10898 ( .B1(n10543), .B2(n10073), .A(n10012), .ZN(n10013) );
  OAI21_X1 U10899 ( .B1(n10014), .B2(n10064), .A(n10013), .ZN(P1_U3228) );
  INV_X1 U10900 ( .A(n9929), .ZN(n10017) );
  NOR3_X1 U10901 ( .A1(n10017), .A2(n10016), .A3(n10015), .ZN(n10020) );
  INV_X1 U10902 ( .A(n10018), .ZN(n10019) );
  OAI21_X1 U10903 ( .B1(n10020), .B2(n10019), .A(n10081), .ZN(n10024) );
  AOI22_X1 U10904 ( .A1(n10087), .A2(n10351), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10023) );
  AOI22_X1 U10905 ( .A1(n10072), .A2(n10380), .B1(n10071), .B2(n10345), .ZN(
        n10022) );
  NAND2_X1 U10906 ( .A1(n10514), .A2(n10073), .ZN(n10021) );
  NAND4_X1 U10907 ( .A1(n10024), .A2(n10023), .A3(n10022), .A4(n10021), .ZN(
        P1_U3229) );
  XOR2_X1 U10908 ( .A(n10026), .B(n10025), .Z(n10034) );
  INV_X1 U10909 ( .A(n10405), .ZN(n10031) );
  OR2_X1 U10910 ( .A1(n10263), .A2(n10462), .ZN(n10028) );
  OR2_X1 U10911 ( .A1(n10433), .A2(n10464), .ZN(n10027) );
  NAND2_X1 U10912 ( .A1(n10028), .A2(n10027), .ZN(n10411) );
  AOI22_X1 U10913 ( .A1(n10411), .A2(n10029), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10030) );
  OAI21_X1 U10914 ( .B1(n10031), .B2(n10084), .A(n10030), .ZN(n10032) );
  AOI21_X1 U10915 ( .B1(n10537), .B2(n10073), .A(n10032), .ZN(n10033) );
  OAI21_X1 U10916 ( .B1(n10034), .B2(n10064), .A(n10033), .ZN(P1_U3233) );
  AND2_X1 U10917 ( .A1(n9803), .A2(n10035), .ZN(n10038) );
  OAI211_X1 U10918 ( .C1(n10038), .C2(n10037), .A(n10081), .B(n10036), .ZN(
        n10046) );
  INV_X1 U10919 ( .A(n10039), .ZN(n10042) );
  OAI21_X1 U10920 ( .B1(n10042), .B2(n10041), .A(n10040), .ZN(n10043) );
  AOI21_X1 U10921 ( .B1(n10044), .B2(n10071), .A(n10043), .ZN(n10045) );
  OAI211_X1 U10922 ( .C1(n10968), .C2(n10090), .A(n10046), .B(n10045), .ZN(
        P1_U3234) );
  NAND2_X1 U10923 ( .A1(n10048), .A2(n10047), .ZN(n10050) );
  XNOR2_X1 U10924 ( .A(n10050), .B(n10049), .ZN(n10056) );
  OAI22_X1 U10925 ( .A1(n10061), .A2(n10267), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10051), .ZN(n10054) );
  INV_X1 U10926 ( .A(n10374), .ZN(n10052) );
  OAI22_X1 U10927 ( .A1(n10085), .A2(n10263), .B1(n10084), .B2(n10052), .ZN(
        n10053) );
  AOI211_X1 U10928 ( .C1(n10525), .C2(n10073), .A(n10054), .B(n10053), .ZN(
        n10055) );
  OAI21_X1 U10929 ( .B1(n10056), .B2(n10064), .A(n10055), .ZN(P1_U3235) );
  AOI21_X1 U10930 ( .B1(n10059), .B2(n10058), .A(n10057), .ZN(n10065) );
  AOI22_X1 U10931 ( .A1(n10072), .A2(n10258), .B1(n10071), .B2(n10439), .ZN(
        n10060) );
  NAND2_X1 U10932 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10201)
         );
  OAI211_X1 U10933 ( .C1(n10061), .C2(n10433), .A(n10060), .B(n10201), .ZN(
        n10062) );
  AOI21_X1 U10934 ( .B1(n10260), .B2(n10073), .A(n10062), .ZN(n10063) );
  OAI21_X1 U10935 ( .B1(n10065), .B2(n10064), .A(n10063), .ZN(P1_U3238) );
  INV_X1 U10936 ( .A(n9982), .ZN(n10068) );
  OAI21_X1 U10937 ( .B1(n10068), .B2(n10067), .A(n10066), .ZN(n10070) );
  NAND3_X1 U10938 ( .A1(n10070), .A2(n10081), .A3(n10069), .ZN(n10077) );
  INV_X1 U10939 ( .A(n10319), .ZN(n10270) );
  AOI22_X1 U10940 ( .A1(n10087), .A2(n10270), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10076) );
  AOI22_X1 U10941 ( .A1(n10072), .A2(n10351), .B1(n10071), .B2(n10323), .ZN(
        n10075) );
  NAND2_X1 U10942 ( .A1(n10506), .A2(n10073), .ZN(n10074) );
  NAND4_X1 U10943 ( .A1(n10077), .A2(n10076), .A3(n10075), .A4(n10074), .ZN(
        P1_U3240) );
  INV_X1 U10944 ( .A(n10556), .ZN(n10996) );
  OAI21_X1 U10945 ( .B1(n10080), .B2(n10079), .A(n10078), .ZN(n10082) );
  NAND2_X1 U10946 ( .A1(n10082), .A2(n10081), .ZN(n10089) );
  AND2_X1 U10947 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10150) );
  INV_X1 U10948 ( .A(n10993), .ZN(n10083) );
  OAI22_X1 U10949 ( .A1(n10085), .A2(n10257), .B1(n10084), .B2(n10083), .ZN(
        n10086) );
  AOI211_X1 U10950 ( .C1(n10087), .C2(n10553), .A(n10150), .B(n10086), .ZN(
        n10088) );
  OAI211_X1 U10951 ( .C1(n10996), .C2(n10090), .A(n10089), .B(n10088), .ZN(
        P1_U3241) );
  MUX2_X1 U10952 ( .A(n10091), .B(P1_DATAO_REG_31__SCAN_IN), .S(n10104), .Z(
        P1_U3585) );
  MUX2_X1 U10953 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n10092), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10954 ( .A(n10271), .B(P1_DATAO_REG_28__SCAN_IN), .S(n10104), .Z(
        P1_U3582) );
  MUX2_X1 U10955 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n10270), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10956 ( .A(n10351), .B(P1_DATAO_REG_25__SCAN_IN), .S(n10104), .Z(
        P1_U3579) );
  MUX2_X1 U10957 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n10363), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10958 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n10389), .S(P1_U3973), .Z(
        P1_U3576) );
  INV_X1 U10959 ( .A(n10263), .ZN(n10381) );
  MUX2_X1 U10960 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n10381), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10961 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n5699), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10962 ( .A(n10417), .B(P1_DATAO_REG_18__SCAN_IN), .S(n10104), .Z(
        P1_U3572) );
  MUX2_X1 U10963 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n10258), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10964 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n10553), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10965 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n5693), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10966 ( .A(n10551), .B(P1_DATAO_REG_14__SCAN_IN), .S(n10104), .Z(
        P1_U3568) );
  MUX2_X1 U10967 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n10093), .S(P1_U3973), .Z(
        P1_U3567) );
  INV_X1 U10968 ( .A(n10094), .ZN(n10095) );
  MUX2_X1 U10969 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n10095), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10970 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n10096), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10971 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n10097), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10972 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n10098), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10973 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n10099), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10974 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n10100), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10975 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n10101), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10976 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n10102), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10977 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n10103), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10978 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n7812), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10979 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n7077), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10980 ( .A(n7973), .B(P1_DATAO_REG_0__SCAN_IN), .S(n10104), .Z(
        P1_U3554) );
  INV_X1 U10981 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10108) );
  NAND2_X1 U10982 ( .A1(n10770), .A2(n10105), .ZN(n10107) );
  NAND2_X1 U10983 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n10106)
         );
  OAI211_X1 U10984 ( .C1(n10108), .C2(n10203), .A(n10107), .B(n10106), .ZN(
        n10109) );
  INV_X1 U10985 ( .A(n10109), .ZN(n10118) );
  OAI211_X1 U10986 ( .C1(n10112), .C2(n10111), .A(n10222), .B(n10110), .ZN(
        n10117) );
  OAI211_X1 U10987 ( .C1(n10115), .C2(n10114), .A(n10147), .B(n10113), .ZN(
        n10116) );
  NAND3_X1 U10988 ( .A1(n10118), .A2(n10117), .A3(n10116), .ZN(P1_U3253) );
  INV_X1 U10989 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10121) );
  NAND2_X1 U10990 ( .A1(n10770), .A2(n10143), .ZN(n10120) );
  OAI211_X1 U10991 ( .C1(n10121), .C2(n10203), .A(n10120), .B(n10119), .ZN(
        n10122) );
  INV_X1 U10992 ( .A(n10122), .ZN(n10136) );
  XNOR2_X1 U10993 ( .A(n10131), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n10126) );
  OAI211_X1 U10994 ( .C1(n10126), .C2(n10125), .A(n10222), .B(n10138), .ZN(
        n10135) );
  INV_X1 U10995 ( .A(n10127), .ZN(n10128) );
  OAI21_X1 U10996 ( .B1(n10129), .B2(n10971), .A(n10128), .ZN(n10133) );
  NAND2_X1 U10997 ( .A1(n10131), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n10130) );
  OAI21_X1 U10998 ( .B1(n10131), .B2(P1_REG1_REG_14__SCAN_IN), .A(n10130), 
        .ZN(n10132) );
  NAND2_X1 U10999 ( .A1(n10132), .A2(n10133), .ZN(n10145) );
  OAI211_X1 U11000 ( .C1(n10133), .C2(n10132), .A(n10147), .B(n10145), .ZN(
        n10134) );
  NAND3_X1 U11001 ( .A1(n10136), .A2(n10135), .A3(n10134), .ZN(P1_U3257) );
  INV_X1 U11002 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10142) );
  NAND2_X1 U11003 ( .A1(n10143), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10137) );
  NAND2_X1 U11004 ( .A1(n10138), .A2(n10137), .ZN(n10140) );
  INV_X1 U11005 ( .A(n10169), .ZN(n10139) );
  OAI21_X1 U11006 ( .B1(n10158), .B2(n10140), .A(n10139), .ZN(n10141) );
  NOR2_X1 U11007 ( .A1(n10142), .A2(n10141), .ZN(n10168) );
  AOI211_X1 U11008 ( .C1(n10142), .C2(n10141), .A(n10168), .B(n10763), .ZN(
        n10156) );
  NAND2_X1 U11009 ( .A1(n10143), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n10144) );
  NAND2_X1 U11010 ( .A1(n10145), .A2(n10144), .ZN(n10159) );
  INV_X1 U11011 ( .A(n10158), .ZN(n10146) );
  XNOR2_X1 U11012 ( .A(n10159), .B(n10146), .ZN(n10148) );
  NAND2_X1 U11013 ( .A1(n10148), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n10161) );
  OAI211_X1 U11014 ( .C1(n10148), .C2(P1_REG1_REG_15__SCAN_IN), .A(n10147), 
        .B(n10161), .ZN(n10149) );
  INV_X1 U11015 ( .A(n10149), .ZN(n10155) );
  INV_X1 U11016 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10153) );
  NAND2_X1 U11017 ( .A1(n10770), .A2(n10158), .ZN(n10152) );
  INV_X1 U11018 ( .A(n10150), .ZN(n10151) );
  OAI211_X1 U11019 ( .C1(n10153), .C2(n10203), .A(n10152), .B(n10151), .ZN(
        n10154) );
  OR3_X1 U11020 ( .A1(n10156), .A2(n10155), .A3(n10154), .ZN(P1_U3258) );
  OR2_X1 U11021 ( .A1(n10182), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n10175) );
  NAND2_X1 U11022 ( .A1(n10182), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n10157) );
  NAND2_X1 U11023 ( .A1(n10175), .A2(n10157), .ZN(n10164) );
  NAND2_X1 U11024 ( .A1(n10159), .A2(n10158), .ZN(n10160) );
  NAND2_X1 U11025 ( .A1(n10161), .A2(n10160), .ZN(n10163) );
  INV_X1 U11026 ( .A(n10176), .ZN(n10162) );
  AOI21_X1 U11027 ( .B1(n10164), .B2(n10163), .A(n10162), .ZN(n10172) );
  NOR2_X1 U11028 ( .A1(n10203), .A2(n10165), .ZN(n10166) );
  AOI211_X1 U11029 ( .C1(n10182), .C2(n10770), .A(n10167), .B(n10166), .ZN(
        n10171) );
  OAI211_X1 U11030 ( .C1(n5188), .C2(n5419), .A(n10222), .B(n10181), .ZN(
        n10170) );
  OAI211_X1 U11031 ( .C1(n10172), .C2(n10759), .A(n10171), .B(n10170), .ZN(
        P1_U3259) );
  OR2_X1 U11032 ( .A1(n10198), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n10174) );
  NAND2_X1 U11033 ( .A1(n10198), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n10173) );
  AND2_X1 U11034 ( .A1(n10174), .A2(n10173), .ZN(n10178) );
  NAND2_X1 U11035 ( .A1(n10176), .A2(n10175), .ZN(n10177) );
  NAND2_X1 U11036 ( .A1(n10177), .A2(n10178), .ZN(n10197) );
  OAI21_X1 U11037 ( .B1(n10178), .B2(n10177), .A(n10197), .ZN(n10179) );
  INV_X1 U11038 ( .A(n10179), .ZN(n10191) );
  NOR2_X1 U11039 ( .A1(n10198), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n10180) );
  AOI21_X1 U11040 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n10198), .A(n10180), 
        .ZN(n10184) );
  NAND2_X1 U11041 ( .A1(n10184), .A2(n10183), .ZN(n10192) );
  OAI21_X1 U11042 ( .B1(n10184), .B2(n10183), .A(n10192), .ZN(n10189) );
  INV_X1 U11043 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10187) );
  NAND2_X1 U11044 ( .A1(n10770), .A2(n10198), .ZN(n10186) );
  OAI211_X1 U11045 ( .C1(n10187), .C2(n10203), .A(n10186), .B(n10185), .ZN(
        n10188) );
  AOI21_X1 U11046 ( .B1(n10222), .B2(n10189), .A(n10188), .ZN(n10190) );
  OAI21_X1 U11047 ( .B1(n10191), .B2(n10759), .A(n10190), .ZN(P1_U3260) );
  OAI21_X1 U11048 ( .B1(n10198), .B2(P1_REG2_REG_17__SCAN_IN), .A(n10192), 
        .ZN(n10195) );
  NAND2_X1 U11049 ( .A1(n10209), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n10213) );
  OAI21_X1 U11050 ( .B1(n10209), .B2(P1_REG2_REG_18__SCAN_IN), .A(n10213), 
        .ZN(n10194) );
  OR2_X1 U11051 ( .A1(n10194), .A2(n10195), .ZN(n10214) );
  INV_X1 U11052 ( .A(n10214), .ZN(n10193) );
  AOI211_X1 U11053 ( .C1(n10195), .C2(n10194), .A(n10193), .B(n10763), .ZN(
        n10207) );
  INV_X1 U11054 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n11024) );
  NOR2_X1 U11055 ( .A1(n10209), .A2(n11024), .ZN(n10196) );
  AOI21_X1 U11056 ( .B1(n10209), .B2(n11024), .A(n10196), .ZN(n10200) );
  OAI21_X1 U11057 ( .B1(n10198), .B2(P1_REG1_REG_17__SCAN_IN), .A(n10197), 
        .ZN(n10199) );
  NOR2_X1 U11058 ( .A1(n10199), .A2(n10200), .ZN(n10208) );
  AOI211_X1 U11059 ( .C1(n10200), .C2(n10199), .A(n10208), .B(n10759), .ZN(
        n10206) );
  INV_X1 U11060 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10204) );
  NAND2_X1 U11061 ( .A1(n10770), .A2(n10209), .ZN(n10202) );
  OAI211_X1 U11062 ( .C1(n10204), .C2(n10203), .A(n10202), .B(n10201), .ZN(
        n10205) );
  OR3_X1 U11063 ( .A1(n10207), .A2(n10206), .A3(n10205), .ZN(P1_U3261) );
  INV_X1 U11064 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n11036) );
  MUX2_X1 U11065 ( .A(n11036), .B(P1_REG1_REG_19__SCAN_IN), .S(n10219), .Z(
        n10211) );
  AOI21_X1 U11066 ( .B1(n10209), .B2(P1_REG1_REG_18__SCAN_IN), .A(n10208), 
        .ZN(n10210) );
  XOR2_X1 U11067 ( .A(n10211), .B(n10210), .Z(n10225) );
  INV_X1 U11068 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10212) );
  MUX2_X1 U11069 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n10212), .S(n10219), .Z(
        n10216) );
  NAND2_X1 U11070 ( .A1(n10214), .A2(n10213), .ZN(n10215) );
  XNOR2_X1 U11071 ( .A(n10216), .B(n10215), .ZN(n10223) );
  NAND2_X1 U11072 ( .A1(n10756), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n10217) );
  OAI211_X1 U11073 ( .C1(n10220), .C2(n10219), .A(n10218), .B(n10217), .ZN(
        n10221) );
  AOI21_X1 U11074 ( .B1(n10223), .B2(n10222), .A(n10221), .ZN(n10224) );
  OAI21_X1 U11075 ( .B1(n10225), .B2(n10759), .A(n10224), .ZN(P1_U3262) );
  NAND2_X1 U11076 ( .A1(n10452), .A2(n11020), .ZN(n10438) );
  NOR2_X1 U11077 ( .A1(n10438), .A2(n10428), .ZN(n10402) );
  NAND2_X1 U11078 ( .A1(n10402), .A2(n10407), .ZN(n10403) );
  INV_X1 U11079 ( .A(n10514), .ZN(n10347) );
  NAND2_X1 U11080 ( .A1(n10330), .A2(n10326), .ZN(n10320) );
  XNOR2_X1 U11081 ( .A(n10484), .B(n5109), .ZN(n10227) );
  NAND2_X1 U11082 ( .A1(n10227), .A2(n10949), .ZN(n10483) );
  AND2_X1 U11083 ( .A1(n10228), .A2(P1_B_REG_SCAN_IN), .ZN(n10229) );
  OR2_X1 U11084 ( .A1(n10462), .A2(n10229), .ZN(n10249) );
  OR2_X1 U11085 ( .A1(n10230), .A2(n10249), .ZN(n10485) );
  NOR2_X1 U11086 ( .A1(n10485), .A2(n11005), .ZN(n10234) );
  NOR2_X1 U11087 ( .A1(n10484), .A2(n10995), .ZN(n10231) );
  AOI211_X1 U11088 ( .C1(n11005), .C2(P1_REG2_REG_31__SCAN_IN), .A(n10234), 
        .B(n10231), .ZN(n10232) );
  OAI21_X1 U11089 ( .B1(n10477), .B2(n10483), .A(n10232), .ZN(P1_U3263) );
  OAI211_X1 U11090 ( .C1(n10487), .C2(n10275), .A(n10949), .B(n5109), .ZN(
        n10486) );
  NOR2_X1 U11091 ( .A1(n10487), .A2(n10995), .ZN(n10233) );
  AOI211_X1 U11092 ( .C1(n11005), .C2(P1_REG2_REG_30__SCAN_IN), .A(n10234), 
        .B(n10233), .ZN(n10235) );
  OAI21_X1 U11093 ( .B1(n10477), .B2(n10486), .A(n10235), .ZN(P1_U3264) );
  NAND2_X1 U11094 ( .A1(n10409), .A2(n10410), .ZN(n10408) );
  NAND2_X1 U11095 ( .A1(n10408), .A2(n10236), .ZN(n10387) );
  INV_X1 U11096 ( .A(n10391), .ZN(n10388) );
  NAND2_X1 U11097 ( .A1(n10387), .A2(n10388), .ZN(n10386) );
  NAND2_X1 U11098 ( .A1(n10386), .A2(n10237), .ZN(n10378) );
  NAND2_X1 U11099 ( .A1(n10378), .A2(n10379), .ZN(n10377) );
  INV_X1 U11100 ( .A(n10239), .ZN(n10240) );
  INV_X1 U11101 ( .A(n10245), .ZN(n10246) );
  INV_X1 U11102 ( .A(n10273), .ZN(n10248) );
  NOR2_X1 U11103 ( .A1(n10250), .A2(n10249), .ZN(n10251) );
  OAI21_X1 U11104 ( .B1(n10253), .B2(n10941), .A(n10252), .ZN(n10489) );
  INV_X1 U11105 ( .A(n10489), .ZN(n10282) );
  OAI21_X1 U11106 ( .B1(n10255), .B2(n10551), .A(n10254), .ZN(n10256) );
  OAI21_X1 U11107 ( .B1(n10975), .B2(n10257), .A(n10256), .ZN(n10547) );
  AOI21_X2 U11108 ( .B1(n10446), .B2(n10445), .A(n10259), .ZN(n10437) );
  NAND2_X1 U11109 ( .A1(n10260), .A2(n10417), .ZN(n10261) );
  NAND2_X1 U11110 ( .A1(n10420), .A2(n10419), .ZN(n10421) );
  INV_X1 U11111 ( .A(n10428), .ZN(n11032) );
  INV_X1 U11112 ( .A(n10531), .ZN(n10396) );
  NAND2_X1 U11113 ( .A1(n10529), .A2(n5719), .ZN(n10370) );
  NAND2_X1 U11114 ( .A1(n10265), .A2(n10267), .ZN(n10266) );
  NAND2_X1 U11115 ( .A1(n10268), .A2(n5721), .ZN(n10341) );
  NAND2_X1 U11116 ( .A1(n10510), .A2(n10351), .ZN(n10269) );
  AOI22_X2 U11117 ( .A1(n10329), .A2(n10269), .B1(n10318), .B2(n5390), .ZN(
        n10314) );
  NOR2_X1 U11118 ( .A1(n10495), .A2(n10271), .ZN(n10272) );
  OAI22_X1 U11119 ( .A1(n10284), .A2(n10272), .B1(n10306), .B2(n10290), .ZN(
        n10274) );
  XNOR2_X1 U11120 ( .A(n10274), .B(n10273), .ZN(n10488) );
  NAND2_X1 U11121 ( .A1(n10488), .A2(n10961), .ZN(n10281) );
  AOI211_X1 U11122 ( .C1(n10491), .C2(n10285), .A(n10976), .B(n10275), .ZN(
        n10490) );
  INV_X1 U11123 ( .A(n10491), .ZN(n10278) );
  AOI22_X1 U11124 ( .A1(n11005), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n10276), 
        .B2(n10992), .ZN(n10277) );
  OAI21_X1 U11125 ( .B1(n10278), .B2(n10995), .A(n10277), .ZN(n10279) );
  AOI21_X1 U11126 ( .B1(n10490), .B2(n10959), .A(n10279), .ZN(n10280) );
  OAI211_X1 U11127 ( .C1(n10282), .C2(n10955), .A(n10281), .B(n10280), .ZN(
        P1_U3356) );
  XNOR2_X1 U11128 ( .A(n10284), .B(n10283), .ZN(n10498) );
  INV_X1 U11129 ( .A(n10307), .ZN(n10287) );
  INV_X1 U11130 ( .A(n10285), .ZN(n10286) );
  AOI211_X1 U11131 ( .C1(n10495), .C2(n10287), .A(n10976), .B(n10286), .ZN(
        n10494) );
  AOI22_X1 U11132 ( .A1(n11005), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n10288), 
        .B2(n10992), .ZN(n10289) );
  OAI21_X1 U11133 ( .B1(n10290), .B2(n10995), .A(n10289), .ZN(n10296) );
  XNOR2_X1 U11134 ( .A(n10292), .B(n10291), .ZN(n10294) );
  AOI21_X1 U11135 ( .B1(n10294), .B2(n10821), .A(n10293), .ZN(n10497) );
  NOR2_X1 U11136 ( .A1(n10497), .A2(n11005), .ZN(n10295) );
  AOI211_X1 U11137 ( .C1(n10959), .C2(n10494), .A(n10296), .B(n10295), .ZN(
        n10297) );
  OAI21_X1 U11138 ( .B1(n10498), .B2(n10458), .A(n10297), .ZN(P1_U3265) );
  INV_X1 U11139 ( .A(n10298), .ZN(n10299) );
  AOI21_X1 U11140 ( .B1(n5522), .B2(n10300), .A(n10299), .ZN(n10503) );
  AOI21_X1 U11141 ( .B1(n10303), .B2(n10302), .A(n10301), .ZN(n10304) );
  OAI222_X1 U11142 ( .A1(n10462), .A2(n10306), .B1(n10464), .B2(n10305), .C1(
        n10941), .C2(n10304), .ZN(n10499) );
  AOI211_X1 U11143 ( .C1(n10501), .C2(n10320), .A(n10976), .B(n10307), .ZN(
        n10500) );
  NAND2_X1 U11144 ( .A1(n10500), .A2(n10959), .ZN(n10310) );
  AOI22_X1 U11145 ( .A1(n11005), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n10308), 
        .B2(n10992), .ZN(n10309) );
  OAI211_X1 U11146 ( .C1(n5414), .C2(n10995), .A(n10310), .B(n10309), .ZN(
        n10311) );
  AOI21_X1 U11147 ( .B1(n10499), .B2(n10475), .A(n10311), .ZN(n10312) );
  OAI21_X1 U11148 ( .B1(n10503), .B2(n10458), .A(n10312), .ZN(P1_U3266) );
  OAI21_X1 U11149 ( .B1(n10314), .B2(n10315), .A(n10313), .ZN(n10508) );
  XNOR2_X1 U11150 ( .A(n10316), .B(n10315), .ZN(n10317) );
  OAI222_X1 U11151 ( .A1(n10462), .A2(n10319), .B1(n10464), .B2(n10318), .C1(
        n10317), .C2(n10941), .ZN(n10504) );
  INV_X1 U11152 ( .A(n10330), .ZN(n10322) );
  INV_X1 U11153 ( .A(n10320), .ZN(n10321) );
  AOI211_X1 U11154 ( .C1(n10506), .C2(n10322), .A(n10976), .B(n10321), .ZN(
        n10505) );
  NAND2_X1 U11155 ( .A1(n10505), .A2(n10959), .ZN(n10325) );
  AOI22_X1 U11156 ( .A1(n11005), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n10323), 
        .B2(n10992), .ZN(n10324) );
  OAI211_X1 U11157 ( .C1(n10326), .C2(n10995), .A(n10325), .B(n10324), .ZN(
        n10327) );
  AOI21_X1 U11158 ( .B1(n10504), .B2(n10475), .A(n10327), .ZN(n10328) );
  OAI21_X1 U11159 ( .B1(n10508), .B2(n10458), .A(n10328), .ZN(P1_U3267) );
  XNOR2_X1 U11160 ( .A(n10329), .B(n10334), .ZN(n10513) );
  AOI211_X1 U11161 ( .C1(n10510), .C2(n10343), .A(n10976), .B(n10330), .ZN(
        n10509) );
  AOI22_X1 U11162 ( .A1(n11005), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n10331), 
        .B2(n10992), .ZN(n10332) );
  OAI21_X1 U11163 ( .B1(n5390), .B2(n10995), .A(n10332), .ZN(n10339) );
  OAI21_X1 U11164 ( .B1(n10335), .B2(n10334), .A(n10333), .ZN(n10337) );
  AOI21_X1 U11165 ( .B1(n10337), .B2(n10821), .A(n10336), .ZN(n10512) );
  NOR2_X1 U11166 ( .A1(n10512), .A2(n11005), .ZN(n10338) );
  AOI211_X1 U11167 ( .C1(n10509), .C2(n10959), .A(n10339), .B(n10338), .ZN(
        n10340) );
  OAI21_X1 U11168 ( .B1(n10513), .B2(n10458), .A(n10340), .ZN(P1_U3268) );
  XNOR2_X1 U11169 ( .A(n10341), .B(n10342), .ZN(n10518) );
  INV_X1 U11170 ( .A(n10343), .ZN(n10344) );
  AOI21_X1 U11171 ( .B1(n10514), .B2(n5394), .A(n10344), .ZN(n10515) );
  AOI22_X1 U11172 ( .A1(n11005), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n10345), 
        .B2(n10992), .ZN(n10346) );
  OAI21_X1 U11173 ( .B1(n10347), .B2(n10995), .A(n10346), .ZN(n10354) );
  NAND2_X1 U11174 ( .A1(n10360), .A2(n10348), .ZN(n10350) );
  XNOR2_X1 U11175 ( .A(n10350), .B(n10349), .ZN(n10352) );
  AOI222_X1 U11176 ( .A1(n10821), .A2(n10352), .B1(n10351), .B2(n10552), .C1(
        n10380), .C2(n10550), .ZN(n10517) );
  NOR2_X1 U11177 ( .A1(n10517), .A2(n11005), .ZN(n10353) );
  AOI211_X1 U11178 ( .C1(n10515), .C2(n11001), .A(n10354), .B(n10353), .ZN(
        n10355) );
  OAI21_X1 U11179 ( .B1(n10518), .B2(n10458), .A(n10355), .ZN(P1_U3269) );
  XOR2_X1 U11180 ( .A(n10362), .B(n10356), .Z(n10523) );
  AOI211_X1 U11181 ( .C1(n10520), .C2(n10371), .A(n10976), .B(n10357), .ZN(
        n10519) );
  AOI22_X1 U11182 ( .A1(n11005), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n10358), 
        .B2(n10992), .ZN(n10359) );
  OAI21_X1 U11183 ( .B1(n10265), .B2(n10995), .A(n10359), .ZN(n10366) );
  OAI21_X1 U11184 ( .B1(n10362), .B2(n10361), .A(n10360), .ZN(n10364) );
  AOI222_X1 U11185 ( .A1(n10821), .A2(n10364), .B1(n10363), .B2(n10552), .C1(
        n10389), .C2(n10550), .ZN(n10522) );
  NOR2_X1 U11186 ( .A1(n10522), .A2(n10955), .ZN(n10365) );
  AOI211_X1 U11187 ( .C1(n10519), .C2(n10959), .A(n10366), .B(n10365), .ZN(
        n10367) );
  OAI21_X1 U11188 ( .B1(n10523), .B2(n10458), .A(n10367), .ZN(P1_U3270) );
  OAI21_X1 U11189 ( .B1(n10370), .B2(n10369), .A(n10368), .ZN(n10528) );
  INV_X1 U11190 ( .A(n10393), .ZN(n10373) );
  INV_X1 U11191 ( .A(n10371), .ZN(n10372) );
  AOI211_X1 U11192 ( .C1(n10525), .C2(n10373), .A(n10976), .B(n10372), .ZN(
        n10524) );
  AOI22_X1 U11193 ( .A1(n11005), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n10374), 
        .B2(n10992), .ZN(n10375) );
  OAI21_X1 U11194 ( .B1(n10376), .B2(n10995), .A(n10375), .ZN(n10384) );
  OAI21_X1 U11195 ( .B1(n10379), .B2(n10378), .A(n10377), .ZN(n10382) );
  AOI222_X1 U11196 ( .A1(n10821), .A2(n10382), .B1(n10381), .B2(n10550), .C1(
        n10380), .C2(n10552), .ZN(n10527) );
  NOR2_X1 U11197 ( .A1(n10527), .A2(n10955), .ZN(n10383) );
  AOI211_X1 U11198 ( .C1(n10524), .C2(n10959), .A(n10384), .B(n10383), .ZN(
        n10385) );
  OAI21_X1 U11199 ( .B1(n10528), .B2(n10458), .A(n10385), .ZN(P1_U3271) );
  OAI21_X1 U11200 ( .B1(n10388), .B2(n10387), .A(n10386), .ZN(n10390) );
  AOI222_X1 U11201 ( .A1(n10821), .A2(n10390), .B1(n10389), .B2(n10552), .C1(
        n5699), .C2(n10550), .ZN(n10534) );
  OR2_X1 U11202 ( .A1(n10392), .A2(n10391), .ZN(n10530) );
  NAND3_X1 U11203 ( .A1(n10530), .A2(n10529), .A3(n10961), .ZN(n10399) );
  AOI21_X1 U11204 ( .B1(n10531), .B2(n10403), .A(n10393), .ZN(n10532) );
  AOI22_X1 U11205 ( .A1(n11005), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n10394), 
        .B2(n10992), .ZN(n10395) );
  OAI21_X1 U11206 ( .B1(n10396), .B2(n10995), .A(n10395), .ZN(n10397) );
  AOI21_X1 U11207 ( .B1(n10532), .B2(n11001), .A(n10397), .ZN(n10398) );
  OAI211_X1 U11208 ( .C1(n11005), .C2(n10534), .A(n10399), .B(n10398), .ZN(
        P1_U3272) );
  AOI21_X1 U11209 ( .B1(n10410), .B2(n10401), .A(n10400), .ZN(n10540) );
  INV_X1 U11210 ( .A(n10402), .ZN(n10424) );
  INV_X1 U11211 ( .A(n10403), .ZN(n10404) );
  AOI211_X1 U11212 ( .C1(n10537), .C2(n10424), .A(n10976), .B(n10404), .ZN(
        n10536) );
  AOI22_X1 U11213 ( .A1(n11005), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n10405), 
        .B2(n10992), .ZN(n10406) );
  OAI21_X1 U11214 ( .B1(n10407), .B2(n10995), .A(n10406), .ZN(n10414) );
  OAI21_X1 U11215 ( .B1(n10410), .B2(n10409), .A(n10408), .ZN(n10412) );
  AOI21_X1 U11216 ( .B1(n10412), .B2(n10821), .A(n10411), .ZN(n10539) );
  NOR2_X1 U11217 ( .A1(n10539), .A2(n11005), .ZN(n10413) );
  AOI211_X1 U11218 ( .C1(n10536), .C2(n10959), .A(n10414), .B(n10413), .ZN(
        n10415) );
  OAI21_X1 U11219 ( .B1(n10540), .B2(n10458), .A(n10415), .ZN(P1_U3273) );
  XNOR2_X1 U11220 ( .A(n10416), .B(n10419), .ZN(n10418) );
  AOI222_X1 U11221 ( .A1(n10821), .A2(n10418), .B1(n5699), .B2(n10552), .C1(
        n10417), .C2(n10550), .ZN(n11030) );
  NOR2_X1 U11222 ( .A1(n10420), .A2(n10419), .ZN(n11028) );
  INV_X1 U11223 ( .A(n11028), .ZN(n10422) );
  NAND3_X1 U11224 ( .A1(n10422), .A2(n10421), .A3(n10961), .ZN(n10430) );
  OAI22_X1 U11225 ( .A1(n10475), .A2(n10212), .B1(n10423), .B2(n10472), .ZN(
        n10427) );
  INV_X1 U11226 ( .A(n10438), .ZN(n10425) );
  OAI211_X1 U11227 ( .C1(n11032), .C2(n10425), .A(n10424), .B(n10949), .ZN(
        n11029) );
  NOR2_X1 U11228 ( .A1(n11029), .A2(n10477), .ZN(n10426) );
  AOI211_X1 U11229 ( .C1(n10956), .C2(n10428), .A(n10427), .B(n10426), .ZN(
        n10429) );
  OAI211_X1 U11230 ( .C1(n11005), .C2(n11030), .A(n10430), .B(n10429), .ZN(
        P1_U3274) );
  INV_X1 U11231 ( .A(n10436), .ZN(n10431) );
  XNOR2_X1 U11232 ( .A(n10432), .B(n10431), .ZN(n10435) );
  OAI22_X1 U11233 ( .A1(n10463), .A2(n10464), .B1(n10433), .B2(n10462), .ZN(
        n10434) );
  AOI21_X1 U11234 ( .B1(n10435), .B2(n10821), .A(n10434), .ZN(n11019) );
  XNOR2_X1 U11235 ( .A(n10437), .B(n10436), .ZN(n11023) );
  NAND2_X1 U11236 ( .A1(n11023), .A2(n10961), .ZN(n10444) );
  OAI211_X1 U11237 ( .C1(n10452), .C2(n11020), .A(n10438), .B(n10949), .ZN(
        n11018) );
  INV_X1 U11238 ( .A(n11018), .ZN(n10442) );
  AOI22_X1 U11239 ( .A1(n11005), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10439), 
        .B2(n10992), .ZN(n10440) );
  OAI21_X1 U11240 ( .B1(n11020), .B2(n10995), .A(n10440), .ZN(n10441) );
  AOI21_X1 U11241 ( .B1(n10442), .B2(n10959), .A(n10441), .ZN(n10443) );
  OAI211_X1 U11242 ( .C1(n11005), .C2(n11019), .A(n10444), .B(n10443), .ZN(
        P1_U3275) );
  XNOR2_X1 U11243 ( .A(n10446), .B(n10445), .ZN(n10545) );
  XNOR2_X1 U11244 ( .A(n10448), .B(n10447), .ZN(n10449) );
  OAI222_X1 U11245 ( .A1(n10462), .A2(n10451), .B1(n10464), .B2(n10450), .C1(
        n10449), .C2(n10941), .ZN(n10541) );
  AOI211_X1 U11246 ( .C1(n10543), .C2(n10476), .A(n10976), .B(n10452), .ZN(
        n10542) );
  NAND2_X1 U11247 ( .A1(n10542), .A2(n10959), .ZN(n10455) );
  AOI22_X1 U11248 ( .A1(n11005), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10453), 
        .B2(n10992), .ZN(n10454) );
  OAI211_X1 U11249 ( .C1(n5396), .C2(n10995), .A(n10455), .B(n10454), .ZN(
        n10456) );
  AOI21_X1 U11250 ( .B1(n10541), .B2(n10475), .A(n10456), .ZN(n10457) );
  OAI21_X1 U11251 ( .B1(n10545), .B2(n10458), .A(n10457), .ZN(P1_U3276) );
  NAND2_X1 U11252 ( .A1(n10459), .A2(n10469), .ZN(n10460) );
  NAND2_X1 U11253 ( .A1(n10461), .A2(n10460), .ZN(n10467) );
  OAI22_X1 U11254 ( .A1(n10465), .A2(n10464), .B1(n10463), .B2(n10462), .ZN(
        n10466) );
  AOI21_X1 U11255 ( .B1(n10467), .B2(n10821), .A(n10466), .ZN(n11007) );
  OAI21_X1 U11256 ( .B1(n10470), .B2(n10469), .A(n10468), .ZN(n10471) );
  INV_X1 U11257 ( .A(n10471), .ZN(n11010) );
  NAND2_X1 U11258 ( .A1(n11010), .A2(n10961), .ZN(n10482) );
  INV_X1 U11259 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10474) );
  OAI22_X1 U11260 ( .A1(n10475), .A2(n10474), .B1(n10473), .B2(n10472), .ZN(
        n10479) );
  OAI211_X1 U11261 ( .C1(n5168), .C2(n11008), .A(n10476), .B(n10949), .ZN(
        n11006) );
  NOR2_X1 U11262 ( .A1(n11006), .A2(n10477), .ZN(n10478) );
  AOI211_X1 U11263 ( .C1(n10956), .C2(n10480), .A(n10479), .B(n10478), .ZN(
        n10481) );
  OAI211_X1 U11264 ( .C1(n11005), .C2(n11007), .A(n10482), .B(n10481), .ZN(
        P1_U3277) );
  OAI211_X1 U11265 ( .C1(n10484), .C2(n11031), .A(n10483), .B(n10485), .ZN(
        n10559) );
  MUX2_X1 U11266 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10559), .S(n11037), .Z(
        P1_U3553) );
  OAI211_X1 U11267 ( .C1(n10487), .C2(n11031), .A(n10486), .B(n10485), .ZN(
        n10560) );
  MUX2_X1 U11268 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10560), .S(n11037), .Z(
        P1_U3552) );
  NAND2_X1 U11269 ( .A1(n10488), .A2(n11022), .ZN(n10493) );
  AOI211_X2 U11270 ( .C1(n10557), .C2(n10491), .A(n10490), .B(n10489), .ZN(
        n10492) );
  NAND2_X1 U11271 ( .A1(n10493), .A2(n10492), .ZN(n10561) );
  MUX2_X1 U11272 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10561), .S(n11037), .Z(
        P1_U3551) );
  AOI21_X1 U11273 ( .B1(n10557), .B2(n10495), .A(n10494), .ZN(n10496) );
  OAI211_X1 U11274 ( .C1(n10498), .C2(n11027), .A(n10497), .B(n10496), .ZN(
        n10562) );
  MUX2_X1 U11275 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10562), .S(n11037), .Z(
        P1_U3550) );
  AOI211_X1 U11276 ( .C1(n10557), .C2(n10501), .A(n10500), .B(n10499), .ZN(
        n10502) );
  OAI21_X1 U11277 ( .B1(n10503), .B2(n11027), .A(n10502), .ZN(n10563) );
  MUX2_X1 U11278 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10563), .S(n11037), .Z(
        P1_U3549) );
  AOI211_X1 U11279 ( .C1(n10557), .C2(n10506), .A(n10505), .B(n10504), .ZN(
        n10507) );
  OAI21_X1 U11280 ( .B1(n10508), .B2(n11027), .A(n10507), .ZN(n10564) );
  MUX2_X1 U11281 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10564), .S(n11037), .Z(
        P1_U3548) );
  AOI21_X1 U11282 ( .B1(n10557), .B2(n10510), .A(n10509), .ZN(n10511) );
  OAI211_X1 U11283 ( .C1(n10513), .C2(n11027), .A(n10512), .B(n10511), .ZN(
        n10565) );
  MUX2_X1 U11284 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10565), .S(n11037), .Z(
        P1_U3547) );
  AOI22_X1 U11285 ( .A1(n10515), .A2(n10949), .B1(n10557), .B2(n10514), .ZN(
        n10516) );
  OAI211_X1 U11286 ( .C1(n10518), .C2(n11027), .A(n10517), .B(n10516), .ZN(
        n10566) );
  MUX2_X1 U11287 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10566), .S(n11037), .Z(
        P1_U3546) );
  AOI21_X1 U11288 ( .B1(n10557), .B2(n10520), .A(n10519), .ZN(n10521) );
  OAI211_X1 U11289 ( .C1(n10523), .C2(n11027), .A(n10522), .B(n10521), .ZN(
        n10567) );
  MUX2_X1 U11290 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10567), .S(n11037), .Z(
        P1_U3545) );
  AOI21_X1 U11291 ( .B1(n10557), .B2(n10525), .A(n10524), .ZN(n10526) );
  OAI211_X1 U11292 ( .C1(n10528), .C2(n11027), .A(n10527), .B(n10526), .ZN(
        n10568) );
  MUX2_X1 U11293 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10568), .S(n11037), .Z(
        P1_U3544) );
  NAND3_X1 U11294 ( .A1(n10530), .A2(n10529), .A3(n11022), .ZN(n10535) );
  AOI22_X1 U11295 ( .A1(n10532), .A2(n10949), .B1(n10557), .B2(n10531), .ZN(
        n10533) );
  NAND3_X1 U11296 ( .A1(n10535), .A2(n10534), .A3(n10533), .ZN(n10569) );
  MUX2_X1 U11297 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10569), .S(n11037), .Z(
        P1_U3543) );
  AOI21_X1 U11298 ( .B1(n10557), .B2(n10537), .A(n10536), .ZN(n10538) );
  OAI211_X1 U11299 ( .C1(n10540), .C2(n11027), .A(n10539), .B(n10538), .ZN(
        n10570) );
  MUX2_X1 U11300 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10570), .S(n11037), .Z(
        P1_U3542) );
  AOI211_X1 U11301 ( .C1(n10557), .C2(n10543), .A(n10542), .B(n10541), .ZN(
        n10544) );
  OAI21_X1 U11302 ( .B1(n10545), .B2(n11027), .A(n10544), .ZN(n10571) );
  MUX2_X1 U11303 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10571), .S(n11037), .Z(
        P1_U3539) );
  AOI21_X1 U11304 ( .B1(n10548), .B2(n10547), .A(n10546), .ZN(n10998) );
  XNOR2_X1 U11305 ( .A(n10549), .B(n10548), .ZN(n10554) );
  AOI222_X1 U11306 ( .A1(n10821), .A2(n10554), .B1(n10553), .B2(n10552), .C1(
        n10551), .C2(n10550), .ZN(n10988) );
  AOI21_X1 U11307 ( .B1(n10556), .B2(n10555), .A(n5168), .ZN(n11002) );
  AOI22_X1 U11308 ( .A1(n11002), .A2(n10949), .B1(n10557), .B2(n10556), .ZN(
        n10558) );
  OAI211_X1 U11309 ( .C1(n10998), .C2(n11027), .A(n10988), .B(n10558), .ZN(
        n10572) );
  MUX2_X1 U11310 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10572), .S(n11037), .Z(
        P1_U3537) );
  MUX2_X1 U11311 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10559), .S(n11041), .Z(
        P1_U3521) );
  MUX2_X1 U11312 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10560), .S(n11041), .Z(
        P1_U3520) );
  MUX2_X1 U11313 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10561), .S(n11041), .Z(
        P1_U3519) );
  MUX2_X1 U11314 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10562), .S(n11041), .Z(
        P1_U3518) );
  MUX2_X1 U11315 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10563), .S(n11041), .Z(
        P1_U3517) );
  MUX2_X1 U11316 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10564), .S(n11041), .Z(
        P1_U3516) );
  MUX2_X1 U11317 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10565), .S(n11041), .Z(
        P1_U3515) );
  MUX2_X1 U11318 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10566), .S(n11041), .Z(
        P1_U3514) );
  MUX2_X1 U11319 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10567), .S(n11041), .Z(
        P1_U3513) );
  MUX2_X1 U11320 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10568), .S(n11041), .Z(
        P1_U3512) );
  MUX2_X1 U11321 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10569), .S(n11041), .Z(
        P1_U3511) );
  MUX2_X1 U11322 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10570), .S(n11041), .Z(
        P1_U3510) );
  MUX2_X1 U11323 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10571), .S(n11041), .Z(
        P1_U3504) );
  MUX2_X1 U11324 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10572), .S(n11041), .Z(
        P1_U3498) );
  MUX2_X1 U11325 ( .A(n10575), .B(P1_D_REG_1__SCAN_IN), .S(n10590), .Z(
        P1_U3440) );
  MUX2_X1 U11326 ( .A(n10576), .B(P1_D_REG_0__SCAN_IN), .S(n10590), .Z(
        P1_U3439) );
  INV_X1 U11327 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10577) );
  NAND3_X1 U11328 ( .A1(n10577), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n10579) );
  OAI22_X1 U11329 ( .A1(n10580), .A2(n10579), .B1(n10578), .B2(n8793), .ZN(
        n10581) );
  AOI21_X1 U11330 ( .B1(n7309), .B2(n10582), .A(n10581), .ZN(n10583) );
  INV_X1 U11331 ( .A(n10583), .ZN(P1_U3324) );
  OAI222_X1 U11332 ( .A1(P1_U3086), .A2(n10584), .B1(n8791), .B2(n10586), .C1(
        n10585), .C2(n8793), .ZN(P1_U3325) );
  MUX2_X1 U11333 ( .A(n10587), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U11334 ( .A1(n10590), .A2(P1_D_REG_2__SCAN_IN), .ZN(P1_U3323) );
  AND2_X1 U11335 ( .A1(n10590), .A2(P1_D_REG_3__SCAN_IN), .ZN(P1_U3322) );
  INV_X1 U11336 ( .A(n10590), .ZN(n10589) );
  NOR2_X1 U11337 ( .A1(n10589), .A2(n10588), .ZN(P1_U3321) );
  AND2_X1 U11338 ( .A1(n10590), .A2(P1_D_REG_5__SCAN_IN), .ZN(P1_U3320) );
  AND2_X1 U11339 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10590), .ZN(P1_U3319) );
  AND2_X1 U11340 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10590), .ZN(P1_U3318) );
  AND2_X1 U11341 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10590), .ZN(P1_U3317) );
  AND2_X1 U11342 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10590), .ZN(P1_U3316) );
  AND2_X1 U11343 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10590), .ZN(P1_U3315) );
  AND2_X1 U11344 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10590), .ZN(P1_U3314) );
  AND2_X1 U11345 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10590), .ZN(P1_U3313) );
  AND2_X1 U11346 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10590), .ZN(P1_U3312) );
  AND2_X1 U11347 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10590), .ZN(P1_U3311) );
  AND2_X1 U11348 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10590), .ZN(P1_U3310) );
  AND2_X1 U11349 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10590), .ZN(P1_U3309) );
  AND2_X1 U11350 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10590), .ZN(P1_U3308) );
  AND2_X1 U11351 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10590), .ZN(P1_U3307) );
  AND2_X1 U11352 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10590), .ZN(P1_U3306) );
  AND2_X1 U11353 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10590), .ZN(P1_U3305) );
  AND2_X1 U11354 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10590), .ZN(P1_U3304) );
  AND2_X1 U11355 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10590), .ZN(P1_U3303) );
  AND2_X1 U11356 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10590), .ZN(P1_U3302) );
  AND2_X1 U11357 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10590), .ZN(P1_U3301) );
  AND2_X1 U11358 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10590), .ZN(P1_U3300) );
  AND2_X1 U11359 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10590), .ZN(P1_U3299) );
  AND2_X1 U11360 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10590), .ZN(P1_U3298) );
  AND2_X1 U11361 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10590), .ZN(P1_U3297) );
  AND2_X1 U11362 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10590), .ZN(P1_U3296) );
  AND2_X1 U11363 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10590), .ZN(P1_U3295) );
  AND2_X1 U11364 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10590), .ZN(P1_U3294) );
  XOR2_X1 U11365 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI222_X1 U11366 ( .A1(n10674), .A2(n10594), .B1(n10674), .B2(n10593), .C1(
        n10592), .C2(n10591), .ZN(ADD_1068_U5) );
  AOI21_X1 U11367 ( .B1(n10597), .B2(n10596), .A(n10595), .ZN(ADD_1068_U54) );
  AOI21_X1 U11368 ( .B1(n10600), .B2(n10599), .A(n10598), .ZN(ADD_1068_U53) );
  OAI21_X1 U11369 ( .B1(n10603), .B2(n10602), .A(n10601), .ZN(ADD_1068_U52) );
  OAI21_X1 U11370 ( .B1(n10606), .B2(n10605), .A(n10604), .ZN(ADD_1068_U51) );
  OAI21_X1 U11371 ( .B1(n10609), .B2(n10608), .A(n10607), .ZN(ADD_1068_U50) );
  OAI21_X1 U11372 ( .B1(n10612), .B2(n10611), .A(n10610), .ZN(ADD_1068_U49) );
  OAI21_X1 U11373 ( .B1(n10615), .B2(n10614), .A(n10613), .ZN(ADD_1068_U48) );
  OAI21_X1 U11374 ( .B1(n10618), .B2(n10617), .A(n10616), .ZN(ADD_1068_U47) );
  OAI21_X1 U11375 ( .B1(n10621), .B2(n10620), .A(n10619), .ZN(ADD_1068_U63) );
  OAI21_X1 U11376 ( .B1(n10624), .B2(n10623), .A(n10622), .ZN(ADD_1068_U62) );
  OAI21_X1 U11377 ( .B1(n10627), .B2(n10626), .A(n10625), .ZN(ADD_1068_U61) );
  OAI21_X1 U11378 ( .B1(n10630), .B2(n10629), .A(n10628), .ZN(ADD_1068_U60) );
  OAI21_X1 U11379 ( .B1(n10633), .B2(n10632), .A(n10631), .ZN(ADD_1068_U59) );
  OAI21_X1 U11380 ( .B1(n10636), .B2(n10635), .A(n10634), .ZN(ADD_1068_U58) );
  OAI21_X1 U11381 ( .B1(n10639), .B2(n10638), .A(n10637), .ZN(ADD_1068_U57) );
  OAI21_X1 U11382 ( .B1(n10642), .B2(n10641), .A(n10640), .ZN(ADD_1068_U56) );
  OAI21_X1 U11383 ( .B1(n10645), .B2(n10644), .A(n10643), .ZN(ADD_1068_U55) );
  AOI22_X1 U11384 ( .A1(n10756), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n10656) );
  NAND2_X1 U11385 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10648) );
  AOI211_X1 U11386 ( .C1(n10648), .C2(n10647), .A(n10646), .B(n10759), .ZN(
        n10653) );
  AOI211_X1 U11387 ( .C1(n10651), .C2(n10650), .A(n10649), .B(n10763), .ZN(
        n10652) );
  AOI211_X1 U11388 ( .C1(n10770), .C2(n10654), .A(n10653), .B(n10652), .ZN(
        n10655) );
  NAND2_X1 U11389 ( .A1(n10656), .A2(n10655), .ZN(P1_U3244) );
  AOI22_X1 U11390 ( .A1(P2_U3893), .A2(n10659), .B1(n10658), .B2(n10657), .ZN(
        P2_U3519) );
  XOR2_X1 U11391 ( .A(n10661), .B(n10660), .Z(n10672) );
  XOR2_X1 U11392 ( .A(n10663), .B(n10662), .Z(n10670) );
  NAND2_X1 U11393 ( .A1(n10722), .A2(n5868), .ZN(n10669) );
  INV_X1 U11394 ( .A(n10717), .ZN(n10667) );
  XNOR2_X1 U11395 ( .A(n10665), .B(n10664), .ZN(n10666) );
  AOI22_X1 U11396 ( .A1(n10667), .A2(n10666), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(P2_U3151), .ZN(n10668) );
  OAI211_X1 U11397 ( .C1(n10724), .C2(n10670), .A(n10669), .B(n10668), .ZN(
        n10671) );
  AOI21_X1 U11398 ( .B1(n10729), .B2(n10672), .A(n10671), .ZN(n10673) );
  OAI21_X1 U11399 ( .B1(n10734), .B2(n10674), .A(n10673), .ZN(P2_U3183) );
  INV_X1 U11400 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10692) );
  AOI21_X1 U11401 ( .B1(n5189), .B2(n10676), .A(n10675), .ZN(n10677) );
  NOR2_X1 U11402 ( .A1(n10717), .A2(n10677), .ZN(n10685) );
  AOI21_X1 U11403 ( .B1(n10680), .B2(n10679), .A(n10678), .ZN(n10683) );
  INV_X1 U11404 ( .A(n10681), .ZN(n10682) );
  OAI21_X1 U11405 ( .B1(n10724), .B2(n10683), .A(n10682), .ZN(n10684) );
  AOI211_X1 U11406 ( .C1(n10722), .C2(n10686), .A(n10685), .B(n10684), .ZN(
        n10691) );
  OAI211_X1 U11407 ( .C1(n10689), .C2(n10688), .A(n10687), .B(n10729), .ZN(
        n10690) );
  OAI211_X1 U11408 ( .C1(n10692), .C2(n10734), .A(n10691), .B(n10690), .ZN(
        P2_U3186) );
  INV_X1 U11409 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10711) );
  AOI21_X1 U11410 ( .B1(n10695), .B2(n10694), .A(n10693), .ZN(n10704) );
  AOI21_X1 U11411 ( .B1(n10698), .B2(n10697), .A(n10696), .ZN(n10699) );
  NOR2_X1 U11412 ( .A1(n10699), .A2(n10724), .ZN(n10700) );
  AOI211_X1 U11413 ( .C1(n10722), .C2(n10702), .A(n10701), .B(n10700), .ZN(
        n10703) );
  OAI21_X1 U11414 ( .B1(n10704), .B2(n10717), .A(n10703), .ZN(n10705) );
  INV_X1 U11415 ( .A(n10705), .ZN(n10710) );
  XOR2_X1 U11416 ( .A(n10707), .B(n10706), .Z(n10708) );
  NAND2_X1 U11417 ( .A1(n10708), .A2(n10729), .ZN(n10709) );
  OAI211_X1 U11418 ( .C1(n10711), .C2(n10734), .A(n10710), .B(n10709), .ZN(
        P2_U3187) );
  INV_X1 U11419 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10735) );
  AOI21_X1 U11420 ( .B1(n10876), .B2(n10713), .A(n10712), .ZN(n10725) );
  AOI21_X1 U11421 ( .B1(n10716), .B2(n10715), .A(n10714), .ZN(n10718) );
  NOR2_X1 U11422 ( .A1(n10718), .A2(n10717), .ZN(n10719) );
  AOI211_X1 U11423 ( .C1(n10722), .C2(n10721), .A(n10720), .B(n10719), .ZN(
        n10723) );
  OAI21_X1 U11424 ( .B1(n10725), .B2(n10724), .A(n10723), .ZN(n10726) );
  INV_X1 U11425 ( .A(n10726), .ZN(n10733) );
  AND2_X1 U11426 ( .A1(n10728), .A2(n10727), .ZN(n10730) );
  OAI21_X1 U11427 ( .B1(n10731), .B2(n10730), .A(n10729), .ZN(n10732) );
  OAI211_X1 U11428 ( .C1(n10735), .C2(n10734), .A(n10733), .B(n10732), .ZN(
        P2_U3189) );
  XOR2_X1 U11429 ( .A(n10736), .B(P1_RD_REG_SCAN_IN), .Z(U126) );
  AOI22_X1 U11430 ( .A1(n10756), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10753) );
  AOI211_X1 U11431 ( .C1(n10739), .C2(n10738), .A(n10737), .B(n10759), .ZN(
        n10744) );
  AOI211_X1 U11432 ( .C1(n10742), .C2(n10741), .A(n10740), .B(n10763), .ZN(
        n10743) );
  AOI211_X1 U11433 ( .C1(n10770), .C2(n10745), .A(n10744), .B(n10743), .ZN(
        n10752) );
  NAND2_X1 U11434 ( .A1(n10746), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10747) );
  XNOR2_X1 U11435 ( .A(n10747), .B(n5427), .ZN(n10748) );
  NAND2_X1 U11436 ( .A1(n10748), .A2(n10750), .ZN(n10749) );
  OAI211_X1 U11437 ( .C1(n10751), .C2(n10750), .A(P1_U3973), .B(n10749), .ZN(
        n10771) );
  NAND3_X1 U11438 ( .A1(n10753), .A2(n10752), .A3(n10771), .ZN(P1_U3245) );
  INV_X1 U11439 ( .A(n10754), .ZN(n10755) );
  AOI21_X1 U11440 ( .B1(n10756), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n10755), .ZN(
        n10773) );
  INV_X1 U11441 ( .A(n10757), .ZN(n10762) );
  INV_X1 U11442 ( .A(n10758), .ZN(n10761) );
  AOI211_X1 U11443 ( .C1(n10762), .C2(n10761), .A(n10760), .B(n10759), .ZN(
        n10768) );
  AOI211_X1 U11444 ( .C1(n10766), .C2(n10765), .A(n10764), .B(n10763), .ZN(
        n10767) );
  AOI211_X1 U11445 ( .C1(n10770), .C2(n10769), .A(n10768), .B(n10767), .ZN(
        n10772) );
  NAND3_X1 U11446 ( .A1(n10773), .A2(n10772), .A3(n10771), .ZN(P1_U3247) );
  OAI211_X1 U11447 ( .C1(n10776), .C2(n11031), .A(n10775), .B(n10774), .ZN(
        n10779) );
  AOI21_X1 U11448 ( .B1(n10848), .B2(n10928), .A(n10777), .ZN(n10778) );
  NOR2_X1 U11449 ( .A1(n10779), .A2(n10778), .ZN(n10781) );
  AOI22_X1 U11450 ( .A1(n11037), .A2(n10781), .B1(n7573), .B2(n11035), .ZN(
        P1_U3523) );
  INV_X1 U11451 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10780) );
  AOI22_X1 U11452 ( .A1(n11041), .A2(n10781), .B1(n10780), .B2(n11038), .ZN(
        P1_U3456) );
  XNOR2_X1 U11453 ( .A(n10783), .B(n10782), .ZN(n10798) );
  INV_X1 U11454 ( .A(n10784), .ZN(n10787) );
  INV_X1 U11455 ( .A(n10785), .ZN(n10786) );
  OAI211_X1 U11456 ( .C1(n7799), .C2(n10787), .A(n10786), .B(n10949), .ZN(
        n10796) );
  OAI21_X1 U11457 ( .B1(n7799), .B2(n11031), .A(n10796), .ZN(n10792) );
  XNOR2_X1 U11458 ( .A(n6745), .B(n10788), .ZN(n10790) );
  AOI21_X1 U11459 ( .B1(n10790), .B2(n10821), .A(n10789), .ZN(n10801) );
  INV_X1 U11460 ( .A(n10801), .ZN(n10791) );
  AOI211_X1 U11461 ( .C1(n11022), .C2(n10798), .A(n10792), .B(n10791), .ZN(
        n10794) );
  AOI22_X1 U11462 ( .A1(n11037), .A2(n10794), .B1(n7575), .B2(n11035), .ZN(
        P1_U3524) );
  INV_X1 U11463 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10793) );
  AOI22_X1 U11464 ( .A1(n11041), .A2(n10794), .B1(n10793), .B2(n11038), .ZN(
        P1_U3459) );
  AOI222_X1 U11465 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n11005), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10992), .C1(n10795), .C2(n10956), .ZN(
        n10800) );
  INV_X1 U11466 ( .A(n10796), .ZN(n10797) );
  AOI22_X1 U11467 ( .A1(n10798), .A2(n10961), .B1(n10797), .B2(n10959), .ZN(
        n10799) );
  OAI211_X1 U11468 ( .C1(n11005), .C2(n10801), .A(n10800), .B(n10799), .ZN(
        P1_U3291) );
  AOI22_X1 U11469 ( .A1(n11017), .A2(n10802), .B1(n6101), .B2(n11015), .ZN(
        P2_U3396) );
  INV_X1 U11470 ( .A(n10928), .ZN(n10979) );
  NAND2_X1 U11471 ( .A1(n10807), .A2(n10979), .ZN(n10804) );
  OAI211_X1 U11472 ( .C1(n7806), .C2(n11031), .A(n10804), .B(n10803), .ZN(
        n10806) );
  AOI211_X1 U11473 ( .C1(n10990), .C2(n10807), .A(n10806), .B(n10805), .ZN(
        n10810) );
  INV_X1 U11474 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U11475 ( .A1(n11037), .A2(n10810), .B1(n10808), .B2(n11035), .ZN(
        P1_U3525) );
  INV_X1 U11476 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U11477 ( .A1(n11041), .A2(n10810), .B1(n10809), .B2(n11038), .ZN(
        P1_U3462) );
  AOI22_X1 U11478 ( .A1(n11017), .A2(n10811), .B1(n6129), .B2(n11015), .ZN(
        P2_U3402) );
  XNOR2_X1 U11479 ( .A(n10812), .B(n10818), .ZN(n10832) );
  INV_X1 U11480 ( .A(n10813), .ZN(n10815) );
  OAI211_X1 U11481 ( .C1(n10815), .C2(n10816), .A(n10949), .B(n10814), .ZN(
        n10830) );
  OAI21_X1 U11482 ( .B1(n10816), .B2(n11031), .A(n10830), .ZN(n10824) );
  XOR2_X1 U11483 ( .A(n10818), .B(n10817), .Z(n10822) );
  INV_X1 U11484 ( .A(n10819), .ZN(n10820) );
  AOI21_X1 U11485 ( .B1(n10822), .B2(n10821), .A(n10820), .ZN(n10835) );
  INV_X1 U11486 ( .A(n10835), .ZN(n10823) );
  AOI211_X1 U11487 ( .C1(n11022), .C2(n10832), .A(n10824), .B(n10823), .ZN(
        n10827) );
  AOI22_X1 U11488 ( .A1(n11037), .A2(n10827), .B1(n10825), .B2(n11035), .ZN(
        P1_U3526) );
  INV_X1 U11489 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10826) );
  AOI22_X1 U11490 ( .A1(n11041), .A2(n10827), .B1(n10826), .B2(n11038), .ZN(
        P1_U3465) );
  AOI222_X1 U11491 ( .A1(n10829), .A2(n10956), .B1(P1_REG2_REG_4__SCAN_IN), 
        .B2(n10955), .C1(n10992), .C2(n10828), .ZN(n10834) );
  INV_X1 U11492 ( .A(n10830), .ZN(n10831) );
  AOI22_X1 U11493 ( .A1(n10832), .A2(n10961), .B1(n10831), .B2(n10959), .ZN(
        n10833) );
  OAI211_X1 U11494 ( .C1(n11005), .C2(n10835), .A(n10834), .B(n10833), .ZN(
        P1_U3289) );
  AOI22_X1 U11495 ( .A1(n11017), .A2(n10836), .B1(n6140), .B2(n11015), .ZN(
        P2_U3405) );
  OAI21_X1 U11496 ( .B1(n10838), .B2(n11031), .A(n10837), .ZN(n10839) );
  AOI21_X1 U11497 ( .B1(n10840), .B2(n11022), .A(n10839), .ZN(n10841) );
  AND2_X1 U11498 ( .A1(n10842), .A2(n10841), .ZN(n10845) );
  INV_X1 U11499 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U11500 ( .A1(n11037), .A2(n10845), .B1(n10843), .B2(n11035), .ZN(
        P1_U3527) );
  INV_X1 U11501 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10844) );
  AOI22_X1 U11502 ( .A1(n11041), .A2(n10845), .B1(n10844), .B2(n11038), .ZN(
        P1_U3468) );
  AOI22_X1 U11503 ( .A1(n11017), .A2(n10846), .B1(n6153), .B2(n11015), .ZN(
        P2_U3408) );
  AOI21_X1 U11504 ( .B1(n10848), .B2(n10928), .A(n10847), .ZN(n10852) );
  OAI211_X1 U11505 ( .C1(n8002), .C2(n11031), .A(n10850), .B(n10849), .ZN(
        n10851) );
  NOR2_X1 U11506 ( .A1(n10852), .A2(n10851), .ZN(n10854) );
  AOI22_X1 U11507 ( .A1(n11037), .A2(n10854), .B1(n7579), .B2(n11035), .ZN(
        P1_U3528) );
  INV_X1 U11508 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U11509 ( .A1(n11041), .A2(n10854), .B1(n10853), .B2(n11038), .ZN(
        P1_U3471) );
  INV_X1 U11510 ( .A(n10855), .ZN(n10861) );
  NOR2_X1 U11511 ( .A1(n10855), .A2(n10928), .ZN(n10860) );
  OAI211_X1 U11512 ( .C1(n10858), .C2(n11031), .A(n10857), .B(n10856), .ZN(
        n10859) );
  AOI211_X1 U11513 ( .C1(n10861), .C2(n10990), .A(n10860), .B(n10859), .ZN(
        n10864) );
  INV_X1 U11514 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U11515 ( .A1(n11037), .A2(n10864), .B1(n10862), .B2(n11035), .ZN(
        P1_U3529) );
  INV_X1 U11516 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10863) );
  AOI22_X1 U11517 ( .A1(n11041), .A2(n10864), .B1(n10863), .B2(n11038), .ZN(
        P1_U3474) );
  INV_X1 U11518 ( .A(n10865), .ZN(n10868) );
  OAI21_X1 U11519 ( .B1(n10868), .B2(n10867), .A(n10866), .ZN(n10873) );
  AOI222_X1 U11520 ( .A1(n10874), .A2(n10873), .B1(n10872), .B2(n10871), .C1(
        n10870), .C2(n10869), .ZN(n10875) );
  OAI21_X1 U11521 ( .B1(n10874), .B2(n10876), .A(n10875), .ZN(P2_U3226) );
  XNOR2_X1 U11522 ( .A(n10877), .B(n10890), .ZN(n10903) );
  INV_X1 U11523 ( .A(n10878), .ZN(n10880) );
  OAI211_X1 U11524 ( .C1(n10880), .C2(n10881), .A(n10949), .B(n10879), .ZN(
        n10900) );
  OAI21_X1 U11525 ( .B1(n10881), .B2(n11031), .A(n10900), .ZN(n10894) );
  NAND2_X1 U11526 ( .A1(n10883), .A2(n10882), .ZN(n10889) );
  INV_X1 U11527 ( .A(n10884), .ZN(n10886) );
  NOR3_X1 U11528 ( .A1(n10887), .A2(n10886), .A3(n10885), .ZN(n10888) );
  AOI211_X1 U11529 ( .C1(n10890), .C2(n10889), .A(n10941), .B(n10888), .ZN(
        n10891) );
  AOI211_X1 U11530 ( .C1(n10990), .C2(n10903), .A(n10892), .B(n10891), .ZN(
        n10906) );
  INV_X1 U11531 ( .A(n10906), .ZN(n10893) );
  AOI211_X1 U11532 ( .C1(n10979), .C2(n10903), .A(n10894), .B(n10893), .ZN(
        n10897) );
  INV_X1 U11533 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U11534 ( .A1(n11037), .A2(n10897), .B1(n10895), .B2(n11035), .ZN(
        P1_U3530) );
  INV_X1 U11535 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10896) );
  AOI22_X1 U11536 ( .A1(n11041), .A2(n10897), .B1(n10896), .B2(n11038), .ZN(
        P1_U3477) );
  AOI222_X1 U11537 ( .A1(n10899), .A2(n10956), .B1(P1_REG2_REG_8__SCAN_IN), 
        .B2(n10955), .C1(n10992), .C2(n10898), .ZN(n10905) );
  INV_X1 U11538 ( .A(n10900), .ZN(n10901) );
  AOI22_X1 U11539 ( .A1(n10903), .A2(n10902), .B1(n10959), .B2(n10901), .ZN(
        n10904) );
  OAI211_X1 U11540 ( .C1(n11005), .C2(n10906), .A(n10905), .B(n10904), .ZN(
        P1_U3285) );
  OAI21_X1 U11541 ( .B1(n10908), .B2(n11031), .A(n10907), .ZN(n10910) );
  AOI211_X1 U11542 ( .C1(n11022), .C2(n10911), .A(n10910), .B(n10909), .ZN(
        n10914) );
  INV_X1 U11543 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U11544 ( .A1(n11037), .A2(n10914), .B1(n10912), .B2(n11035), .ZN(
        P1_U3531) );
  INV_X1 U11545 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10913) );
  AOI22_X1 U11546 ( .A1(n11041), .A2(n10914), .B1(n10913), .B2(n11038), .ZN(
        P1_U3480) );
  OAI211_X1 U11547 ( .C1(n10917), .C2(n11031), .A(n10916), .B(n10915), .ZN(
        n10918) );
  AOI21_X1 U11548 ( .B1(n10919), .B2(n11022), .A(n10918), .ZN(n10922) );
  AOI22_X1 U11549 ( .A1(n11037), .A2(n10922), .B1(n10920), .B2(n11035), .ZN(
        P1_U3532) );
  INV_X1 U11550 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10921) );
  AOI22_X1 U11551 ( .A1(n11041), .A2(n10922), .B1(n10921), .B2(n11038), .ZN(
        P1_U3483) );
  AOI22_X1 U11552 ( .A1(n11017), .A2(n10923), .B1(n6211), .B2(n11015), .ZN(
        P2_U3420) );
  AOI22_X1 U11553 ( .A1(n11017), .A2(n10924), .B1(n6224), .B2(n11015), .ZN(
        P2_U3423) );
  OAI211_X1 U11554 ( .C1(n10927), .C2(n11031), .A(n10926), .B(n10925), .ZN(
        n10931) );
  NOR2_X1 U11555 ( .A1(n10929), .A2(n10928), .ZN(n10930) );
  AOI211_X1 U11556 ( .C1(n10990), .C2(n10932), .A(n10931), .B(n10930), .ZN(
        n10935) );
  AOI22_X1 U11557 ( .A1(n11037), .A2(n10935), .B1(n10933), .B2(n11035), .ZN(
        P1_U3533) );
  INV_X1 U11558 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U11559 ( .A1(n11041), .A2(n10935), .B1(n10934), .B2(n11038), .ZN(
        P1_U3486) );
  AOI22_X1 U11560 ( .A1(n11017), .A2(n10936), .B1(n6235), .B2(n11015), .ZN(
        P2_U3426) );
  XNOR2_X1 U11561 ( .A(n10937), .B(n10938), .ZN(n10962) );
  NOR2_X1 U11562 ( .A1(n10940), .A2(n5526), .ZN(n10942) );
  AOI21_X1 U11563 ( .B1(n10943), .B2(n10942), .A(n10941), .ZN(n10945) );
  AOI21_X1 U11564 ( .B1(n10946), .B2(n10945), .A(n10944), .ZN(n10965) );
  OAI211_X1 U11565 ( .C1(n5406), .C2(n10950), .A(n10949), .B(n10948), .ZN(
        n10958) );
  OAI211_X1 U11566 ( .C1(n10950), .C2(n11031), .A(n10965), .B(n10958), .ZN(
        n10951) );
  AOI21_X1 U11567 ( .B1(n10962), .B2(n11022), .A(n10951), .ZN(n10953) );
  AOI22_X1 U11568 ( .A1(n11037), .A2(n10953), .B1(n8385), .B2(n11035), .ZN(
        P1_U3534) );
  INV_X1 U11569 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10952) );
  AOI22_X1 U11570 ( .A1(n11041), .A2(n10953), .B1(n10952), .B2(n11038), .ZN(
        P1_U3489) );
  AOI222_X1 U11571 ( .A1(n10957), .A2(n10956), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n10955), .C1(n10992), .C2(n10954), .ZN(n10964) );
  INV_X1 U11572 ( .A(n10958), .ZN(n10960) );
  AOI22_X1 U11573 ( .A1(n10962), .A2(n10961), .B1(n10960), .B2(n10959), .ZN(
        n10963) );
  OAI211_X1 U11574 ( .C1(n11005), .C2(n10965), .A(n10964), .B(n10963), .ZN(
        P1_U3281) );
  OAI211_X1 U11575 ( .C1(n10968), .C2(n11031), .A(n10967), .B(n10966), .ZN(
        n10969) );
  AOI21_X1 U11576 ( .B1(n10970), .B2(n11022), .A(n10969), .ZN(n10973) );
  AOI22_X1 U11577 ( .A1(n11037), .A2(n10973), .B1(n10971), .B2(n11035), .ZN(
        P1_U3535) );
  INV_X1 U11578 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10972) );
  AOI22_X1 U11579 ( .A1(n11041), .A2(n10973), .B1(n10972), .B2(n11038), .ZN(
        P1_U3492) );
  AOI22_X1 U11580 ( .A1(n11017), .A2(n10974), .B1(n6248), .B2(n11015), .ZN(
        P2_U3429) );
  OAI22_X1 U11581 ( .A1(n10977), .A2(n10976), .B1(n10975), .B2(n11031), .ZN(
        n10978) );
  AOI21_X1 U11582 ( .B1(n10980), .B2(n10979), .A(n10978), .ZN(n10981) );
  AND2_X1 U11583 ( .A1(n10982), .A2(n10981), .ZN(n10985) );
  INV_X1 U11584 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10983) );
  AOI22_X1 U11585 ( .A1(n11037), .A2(n10985), .B1(n10983), .B2(n11035), .ZN(
        P1_U3536) );
  INV_X1 U11586 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10984) );
  AOI22_X1 U11587 ( .A1(n11041), .A2(n10985), .B1(n10984), .B2(n11038), .ZN(
        P1_U3495) );
  AOI22_X1 U11588 ( .A1(n11017), .A2(n10986), .B1(n6260), .B2(n11015), .ZN(
        P2_U3432) );
  AOI22_X1 U11589 ( .A1(n11017), .A2(n10987), .B1(n6272), .B2(n11015), .ZN(
        P2_U3435) );
  INV_X1 U11590 ( .A(n10998), .ZN(n10991) );
  INV_X1 U11591 ( .A(n10988), .ZN(n10989) );
  AOI21_X1 U11592 ( .B1(n10991), .B2(n10990), .A(n10989), .ZN(n11004) );
  AOI22_X1 U11593 ( .A1(n11005), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n10993), 
        .B2(n10992), .ZN(n10994) );
  OAI21_X1 U11594 ( .B1(n10996), .B2(n10995), .A(n10994), .ZN(n11000) );
  NOR2_X1 U11595 ( .A1(n10998), .A2(n10997), .ZN(n10999) );
  AOI211_X1 U11596 ( .C1(n11002), .C2(n11001), .A(n11000), .B(n10999), .ZN(
        n11003) );
  OAI21_X1 U11597 ( .B1(n11005), .B2(n11004), .A(n11003), .ZN(P1_U3278) );
  OAI211_X1 U11598 ( .C1(n11008), .C2(n11031), .A(n11007), .B(n11006), .ZN(
        n11009) );
  AOI21_X1 U11599 ( .B1(n11010), .B2(n11022), .A(n11009), .ZN(n11013) );
  INV_X1 U11600 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11011) );
  AOI22_X1 U11601 ( .A1(n11037), .A2(n11013), .B1(n11011), .B2(n11035), .ZN(
        P1_U3538) );
  INV_X1 U11602 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n11012) );
  AOI22_X1 U11603 ( .A1(n11041), .A2(n11013), .B1(n11012), .B2(n11038), .ZN(
        P1_U3501) );
  AOI22_X1 U11604 ( .A1(n11017), .A2(n11014), .B1(n6286), .B2(n11015), .ZN(
        P2_U3438) );
  AOI22_X1 U11605 ( .A1(n11017), .A2(n11016), .B1(n6300), .B2(n11015), .ZN(
        P2_U3441) );
  OAI211_X1 U11606 ( .C1(n11020), .C2(n11031), .A(n11019), .B(n11018), .ZN(
        n11021) );
  AOI21_X1 U11607 ( .B1(n11023), .B2(n11022), .A(n11021), .ZN(n11026) );
  AOI22_X1 U11608 ( .A1(n11037), .A2(n11026), .B1(n11024), .B2(n11035), .ZN(
        P1_U3540) );
  INV_X1 U11609 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n11025) );
  AOI22_X1 U11610 ( .A1(n11041), .A2(n11026), .B1(n11025), .B2(n11038), .ZN(
        P1_U3507) );
  NOR2_X1 U11611 ( .A1(n11028), .A2(n11027), .ZN(n11034) );
  OAI211_X1 U11612 ( .C1(n11032), .C2(n11031), .A(n11030), .B(n11029), .ZN(
        n11033) );
  AOI21_X1 U11613 ( .B1(n11034), .B2(n10421), .A(n11033), .ZN(n11040) );
  AOI22_X1 U11614 ( .A1(n11037), .A2(n11040), .B1(n11036), .B2(n11035), .ZN(
        P1_U3541) );
  INV_X1 U11615 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n11039) );
  AOI22_X1 U11616 ( .A1(n11041), .A2(n11040), .B1(n11039), .B2(n11038), .ZN(
        P1_U3509) );
  XNOR2_X1 U11617 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  AND2_X1 U6456 ( .A1(n5207), .A2(n5206), .ZN(n9547) );
endmodule

