

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput63,
         keyinput62, keyinput61, keyinput60, keyinput59, keyinput58,
         keyinput57, keyinput56, keyinput55, keyinput54, keyinput53,
         keyinput52, keyinput51, keyinput50, keyinput49, keyinput48,
         keyinput47, keyinput46, keyinput45, keyinput44, keyinput43,
         keyinput42, keyinput41, keyinput40, keyinput39, keyinput38,
         keyinput37, keyinput36, keyinput35, keyinput34, keyinput33,
         keyinput32, keyinput31, keyinput30, keyinput29, keyinput28,
         keyinput27, keyinput26, keyinput25, keyinput24, keyinput23,
         keyinput22, keyinput21, keyinput20, keyinput19, keyinput18,
         keyinput17, keyinput16, keyinput15, keyinput14, keyinput13,
         keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7,
         keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1,
         keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259;

  AOI211_X1 U7168 ( .C1(n12490), .C2(n12489), .A(n12488), .B(n12487), .ZN(
        n12492) );
  NAND2_X1 U7169 ( .A1(n12561), .A2(n12560), .ZN(n12640) );
  INV_X4 U7170 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7171 ( .A(n12897), .ZN(n13111) );
  OR2_X1 U7172 ( .A1(n10293), .A2(n12227), .ZN(n10319) );
  AND2_X1 U7173 ( .A1(n14132), .A2(n9228), .ZN(n9242) );
  INV_X1 U7174 ( .A(n9326), .ZN(n6649) );
  AND2_X1 U7175 ( .A1(n9343), .A2(n9342), .ZN(n9745) );
  INV_X2 U7176 ( .A(n10055), .ZN(n12548) );
  CLKBUF_X2 U7177 ( .A(n7974), .Z(n9876) );
  CLKBUF_X1 U7178 ( .A(n12273), .Z(n6651) );
  NAND2_X2 U7179 ( .A1(n9843), .A2(n9842), .ZN(n12268) );
  OAI21_X2 U7180 ( .B1(n8834), .B2(n8833), .A(n8832), .ZN(n9028) );
  NAND2_X2 U7181 ( .A1(n9707), .A2(n9706), .ZN(n12259) );
  NAND2_X1 U7182 ( .A1(n8605), .A2(n13574), .ZN(n10313) );
  INV_X1 U7183 ( .A(n6667), .ZN(n12498) );
  NAND2_X1 U7184 ( .A1(n7612), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7611) );
  INV_X1 U7185 ( .A(n12397), .ZN(n12412) );
  INV_X1 U7186 ( .A(n8931), .ZN(n11504) );
  INV_X2 U7187 ( .A(n12399), .ZN(n12393) );
  INV_X2 U7188 ( .A(n12400), .ZN(n11505) );
  OAI211_X2 U7189 ( .C1(n12400), .C2(n8846), .A(n8845), .B(n8844), .ZN(n13916)
         );
  NAND2_X1 U7190 ( .A1(n12489), .A2(n10750), .ZN(n15101) );
  INV_X1 U7191 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8323) );
  NOR2_X1 U7192 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n8165) );
  NOR2_X1 U7193 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n8164) );
  NOR2_X1 U7194 ( .A1(n8214), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n8139) );
  NAND2_X1 U7195 ( .A1(n8137), .A2(n8138), .ZN(n8214) );
  NOR2_X1 U7196 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n8134) );
  AND2_X1 U7197 ( .A1(n11980), .A2(n11979), .ZN(n6456) );
  INV_X1 U7198 ( .A(n12917), .ZN(n12919) );
  NOR2_X1 U7199 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n8133) );
  INV_X1 U7200 ( .A(n11933), .ZN(n12124) );
  INV_X1 U7201 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8366) );
  AND2_X1 U7202 ( .A1(n7681), .A2(n7595), .ZN(n7654) );
  XNOR2_X1 U7203 ( .A(n13916), .B(n13560), .ZN(n12453) );
  INV_X1 U7204 ( .A(n11870), .ZN(n11880) );
  INV_X1 U7205 ( .A(n7750), .ZN(n8005) );
  INV_X1 U7206 ( .A(n9135), .ZN(n7947) );
  AND2_X1 U7207 ( .A1(n11066), .A2(n7231), .ZN(n7230) );
  INV_X1 U7208 ( .A(n9352), .ZN(n11618) );
  NAND2_X1 U7209 ( .A1(n8933), .A2(n8932), .ZN(n15089) );
  OR2_X1 U7210 ( .A1(n10379), .A2(n12399), .ZN(n9707) );
  XNOR2_X1 U7211 ( .A(n6947), .B(n8586), .ZN(n8606) );
  CLKBUF_X3 U7212 ( .A(n9592), .Z(n9593) );
  OR2_X1 U7213 ( .A1(n8715), .A2(n8964), .ZN(n8967) );
  INV_X1 U7214 ( .A(n11874), .ZN(n11879) );
  AND4_X1 U7215 ( .A1(n7695), .A2(n7694), .A3(n7693), .A4(n7692), .ZN(n9780)
         );
  OR2_X1 U7216 ( .A1(n8029), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n8068) );
  NAND2_X1 U7217 ( .A1(n10405), .A2(n10404), .ZN(n14017) );
  BUF_X1 U7218 ( .A(n12488), .Z(n12441) );
  NAND2_X1 U7219 ( .A1(n14196), .A2(n14195), .ZN(n14194) );
  XNOR2_X1 U7220 ( .A(n7353), .B(n6540), .ZN(n14232) );
  CLKBUF_X2 U7221 ( .A(n11435), .Z(n6575) );
  XNOR2_X1 U7222 ( .A(n8178), .B(P1_IR_REG_25__SCAN_IN), .ZN(n14692) );
  NAND3_X1 U7223 ( .A1(n8609), .A2(n8610), .A3(n6961), .ZN(n13561) );
  AOI211_X1 U7224 ( .C1(P2_ADDR_REG_19__SCAN_IN), .C2(n14987), .A(n13577), .B(
        n13576), .ZN(n13578) );
  INV_X1 U7225 ( .A(n15112), .ZN(n15109) );
  NAND4_X1 U7226 ( .A1(n9237), .A2(n9236), .A3(n9235), .A4(n9234), .ZN(n14263)
         );
  AND3_X1 U7227 ( .A1(n6792), .A2(n6626), .A3(n14347), .ZN(n14574) );
  AND4_X1 U7228 ( .A1(n8146), .A2(n8145), .A3(n8144), .A4(n8143), .ZN(n6420)
         );
  XOR2_X1 U7229 ( .A(n9844), .B(n9845), .Z(n6421) );
  NAND2_X1 U7230 ( .A1(n13482), .A2(n13481), .ZN(n13480) );
  AOI21_X2 U7231 ( .B1(n9397), .B2(n9396), .A(n7414), .ZN(n9522) );
  BUF_X4 U7232 ( .A(n7750), .Z(n6422) );
  NAND2_X1 U7233 ( .A1(n9135), .A2(n11907), .ZN(n7750) );
  NAND2_X2 U7234 ( .A1(n7519), .A2(n7518), .ZN(n14863) );
  OAI21_X2 U7235 ( .B1(n10546), .B2(n7259), .A(n7258), .ZN(n10829) );
  AOI21_X2 U7236 ( .B1(n11626), .B2(n13891), .A(n11625), .ZN(n13946) );
  OAI21_X2 U7237 ( .B1(n7146), .B2(n6703), .A(n6701), .ZN(n7814) );
  AOI21_X2 U7238 ( .B1(n9432), .B2(P2_REG1_REG_7__SCAN_IN), .A(n8535), .ZN(
        n15031) );
  XNOR2_X2 U7239 ( .A(n7611), .B(P3_IR_REG_30__SCAN_IN), .ZN(n7618) );
  XNOR2_X2 U7240 ( .A(n11657), .B(n11656), .ZN(n13400) );
  INV_X2 U7241 ( .A(n8975), .ZN(n6423) );
  AND2_X2 U7242 ( .A1(n9248), .A2(n8704), .ZN(n11875) );
  INV_X2 U7243 ( .A(n8975), .ZN(n11825) );
  INV_X4 U7244 ( .A(n11875), .ZN(n8975) );
  NAND2_X2 U7245 ( .A1(n14677), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8690) );
  INV_X1 U7246 ( .A(n13558), .ZN(n8952) );
  NOR2_X2 U7247 ( .A1(n8491), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n8488) );
  AND3_X2 U7248 ( .A1(n9758), .A2(n9746), .A3(n9701), .ZN(n9702) );
  XNOR2_X2 U7249 ( .A(n7661), .B(n7660), .ZN(n9776) );
  AND2_X2 U7250 ( .A1(n12873), .A2(n12874), .ZN(n13188) );
  NAND4_X2 U7251 ( .A1(n8679), .A2(n8678), .A3(n8677), .A4(n8676), .ZN(n13560)
         );
  NAND2_X2 U7252 ( .A1(n14811), .A2(n14810), .ZN(n14822) );
  AOI22_X2 U7253 ( .A1(n14873), .A2(n14874), .B1(n11009), .B2(n11010), .ZN(
        n14811) );
  INV_X2 U7254 ( .A(n13926), .ZN(n12194) );
  XNOR2_X2 U7255 ( .A(n7607), .B(n7606), .ZN(n8045) );
  NOR2_X2 U7256 ( .A1(n14714), .A2(n7508), .ZN(n14719) );
  NOR2_X2 U7257 ( .A1(n14715), .A2(n14716), .ZN(n14714) );
  NOR2_X1 U7258 ( .A1(n10114), .A2(n10115), .ZN(n11003) );
  NAND2_X2 U7259 ( .A1(n8376), .A2(n8375), .ZN(n8463) );
  NOR2_X2 U7260 ( .A1(n10626), .A2(n10625), .ZN(n10628) );
  INV_X1 U7261 ( .A(n15194), .ZN(n10062) );
  XNOR2_X2 U7262 ( .A(n7494), .B(n7493), .ZN(n14711) );
  NAND2_X2 U7263 ( .A1(n15246), .A2(n7492), .ZN(n7494) );
  NOR2_X2 U7264 ( .A1(n8575), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n8573) );
  NOR2_X2 U7265 ( .A1(n8208), .A2(n8705), .ZN(n8230) );
  AOI21_X2 U7266 ( .B1(n10923), .B2(P2_REG1_REG_16__SCAN_IN), .A(n10894), .ZN(
        n10896) );
  XNOR2_X2 U7267 ( .A(n11717), .B(n11716), .ZN(n11695) );
  AOI21_X2 U7268 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(n7510), .A(n14717), .ZN(
        n14844) );
  NOR2_X1 U7269 ( .A1(n14563), .A2(n6946), .ZN(n6945) );
  NAND2_X1 U7270 ( .A1(n13435), .A2(n7411), .ZN(n13482) );
  NAND2_X1 U7271 ( .A1(n13786), .A2(n13791), .ZN(n13788) );
  OAI21_X1 U7272 ( .B1(n14370), .B2(n12153), .A(n6466), .ZN(n14360) );
  NAND2_X1 U7273 ( .A1(n14387), .A2(n14386), .ZN(n14385) );
  NAND2_X1 U7274 ( .A1(n14140), .A2(n11823), .ZN(n14196) );
  NAND2_X1 U7275 ( .A1(n11429), .A2(n11428), .ZN(n14578) );
  NAND2_X1 U7276 ( .A1(n11675), .A2(n7233), .ZN(n13444) );
  AOI21_X1 U7277 ( .B1(n6883), .B2(n6884), .A(n6513), .ZN(n6880) );
  NAND2_X1 U7278 ( .A1(n11329), .A2(n11328), .ZN(n14572) );
  NAND2_X1 U7279 ( .A1(n14165), .A2(n11802), .ZN(n14176) );
  AOI21_X2 U7280 ( .B1(n6886), .B2(n6428), .A(n6512), .ZN(n6885) );
  NAND2_X1 U7281 ( .A1(n7230), .A2(n11067), .ZN(n11104) );
  NAND2_X1 U7282 ( .A1(n11333), .A2(n11332), .ZN(n14586) );
  NAND2_X1 U7283 ( .A1(n14232), .A2(n14231), .ZN(n14230) );
  XNOR2_X1 U7284 ( .A(n11327), .B(n11326), .ZN(n11756) );
  OAI21_X1 U7285 ( .B1(n12944), .B2(n6428), .A(n6467), .ZN(n6879) );
  NAND2_X1 U7286 ( .A1(n11065), .A2(n11064), .ZN(n11066) );
  NAND2_X1 U7287 ( .A1(n11215), .A2(n11214), .ZN(n11785) );
  OAI21_X1 U7288 ( .B1(n12650), .B2(n12648), .A(n13221), .ZN(n12529) );
  NAND2_X1 U7289 ( .A1(n11507), .A2(n11506), .ZN(n13899) );
  NAND2_X1 U7290 ( .A1(n14822), .A2(n11022), .ZN(n14824) );
  NAND2_X1 U7291 ( .A1(n10798), .A2(n7351), .ZN(n11158) );
  NAND2_X1 U7292 ( .A1(n7576), .A2(n6719), .ZN(n7959) );
  OAI22_X1 U7293 ( .A1(n10197), .A2(n10196), .B1(SI_18_), .B2(n10195), .ZN(
        n10201) );
  AND2_X1 U7294 ( .A1(n6720), .A2(n10192), .ZN(n6719) );
  OR2_X1 U7296 ( .A1(n14119), .A2(n11780), .ZN(n12020) );
  NAND2_X1 U7297 ( .A1(n10839), .A2(n10838), .ZN(n14835) );
  NAND2_X1 U7298 ( .A1(n7651), .A2(n7650), .ZN(n7653) );
  NAND2_X1 U7299 ( .A1(n7328), .A2(n7326), .ZN(n10186) );
  NAND2_X1 U7300 ( .A1(n10535), .A2(n10534), .ZN(n14828) );
  XNOR2_X1 U7301 ( .A(n9028), .B(n9027), .ZN(n10830) );
  OAI211_X1 U7302 ( .C1(n14712), .C2(n6737), .A(n6734), .B(n6735), .ZN(n14715)
         );
  NAND2_X1 U7303 ( .A1(n14713), .A2(n15044), .ZN(n14712) );
  NAND2_X1 U7304 ( .A1(n6767), .A2(SI_10_), .ZN(n8631) );
  NAND2_X2 U7306 ( .A1(n6565), .A2(n9484), .ZN(n12245) );
  NAND2_X1 U7307 ( .A1(n8463), .A2(n6435), .ZN(n8464) );
  NAND2_X1 U7308 ( .A1(n6726), .A2(n6728), .ZN(n6731) );
  NAND2_X1 U7309 ( .A1(n8372), .A2(n8371), .ZN(n8376) );
  NAND2_X1 U7310 ( .A1(n8372), .A2(n8355), .ZN(n10098) );
  NAND2_X1 U7311 ( .A1(n9434), .A2(n9433), .ZN(n13414) );
  NAND2_X1 U7312 ( .A1(n9928), .A2(n9927), .ZN(n14096) );
  OR2_X1 U7313 ( .A1(n8354), .A2(n8353), .ZN(n8355) );
  NAND2_X1 U7314 ( .A1(n8354), .A2(n8353), .ZN(n8372) );
  NAND2_X1 U7315 ( .A1(n8350), .A2(n8349), .ZN(n8354) );
  NAND2_X1 U7316 ( .A1(n9388), .A2(n11956), .ZN(n9516) );
  INV_X1 U7317 ( .A(n11964), .ZN(n11966) );
  NAND2_X1 U7318 ( .A1(n9240), .A2(n6795), .ZN(n11964) );
  NAND2_X1 U7319 ( .A1(n10062), .A2(n9778), .ZN(n12777) );
  NAND2_X1 U7320 ( .A1(n6624), .A2(n6864), .ZN(n14135) );
  INV_X1 U7321 ( .A(n9780), .ZN(n15173) );
  OR2_X2 U7322 ( .A1(n9248), .A2(n8187), .ZN(n14266) );
  NAND4_X1 U7323 ( .A1(n7715), .A2(n7714), .A3(n7713), .A4(n7712), .ZN(n15194)
         );
  AOI21_X1 U7324 ( .B1(n6939), .B2(n6438), .A(n6508), .ZN(n6938) );
  CLKBUF_X1 U7325 ( .A(n10313), .Z(n6597) );
  OR2_X1 U7326 ( .A1(n11921), .A2(n8694), .ZN(n8700) );
  OR2_X1 U7327 ( .A1(n9924), .A2(n8969), .ZN(n8970) );
  CLKBUF_X1 U7328 ( .A(n8084), .Z(n11777) );
  AND2_X1 U7329 ( .A1(n9136), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9282) );
  NAND2_X1 U7330 ( .A1(n8176), .A2(n8175), .ZN(n11164) );
  INV_X2 U7331 ( .A(n11793), .ZN(n11881) );
  CLKBUF_X2 U7332 ( .A(n10750), .Z(n6667) );
  BUF_X2 U7333 ( .A(n8996), .Z(n11381) );
  BUF_X2 U7334 ( .A(n11528), .Z(n6638) );
  NAND2_X2 U7335 ( .A1(n9135), .A2(n8968), .ZN(n7749) );
  INV_X1 U7336 ( .A(n8490), .ZN(n10750) );
  OR2_X1 U7337 ( .A1(n11391), .A2(n8204), .ZN(n8971) );
  INV_X1 U7338 ( .A(n14540), .ZN(n11367) );
  NAND2_X1 U7339 ( .A1(n8177), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8178) );
  CLKBUF_X1 U7341 ( .A(n11473), .Z(n6629) );
  XNOR2_X1 U7342 ( .A(n8489), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8490) );
  XNOR2_X1 U7343 ( .A(n8324), .B(n8323), .ZN(n11931) );
  XNOR2_X1 U7344 ( .A(n8703), .B(n8702), .ZN(n12110) );
  XNOR2_X1 U7345 ( .A(n8321), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8784) );
  OR2_X1 U7346 ( .A1(n8488), .A2(n14068), .ZN(n8489) );
  XNOR2_X1 U7347 ( .A(n8492), .B(P2_IR_REG_21__SCAN_IN), .ZN(n12488) );
  XNOR2_X1 U7348 ( .A(n8692), .B(n8691), .ZN(n8693) );
  XNOR2_X1 U7349 ( .A(n8577), .B(n8576), .ZN(n13574) );
  NAND2_X1 U7350 ( .A1(n8591), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8590) );
  NAND2_X1 U7351 ( .A1(n7538), .A2(n7537), .ZN(n7733) );
  CLKBUF_X1 U7352 ( .A(n7654), .Z(n7655) );
  NAND2_X2 U7353 ( .A1(n11907), .A2(P3_U3151), .ZN(n9579) );
  INV_X8 U7354 ( .A(n8968), .ZN(n11907) );
  NAND2_X2 U7355 ( .A1(n8968), .A2(P1_U3086), .ZN(n14694) );
  AND2_X2 U7356 ( .A1(n7313), .A2(n7311), .ZN(n8236) );
  AND4_X1 U7357 ( .A1(n7593), .A2(n7592), .A3(n7807), .A4(n7787), .ZN(n7594)
         );
  AND2_X1 U7358 ( .A1(n8136), .A2(n8135), .ZN(n8261) );
  AND3_X1 U7359 ( .A1(n6823), .A2(n6822), .A3(n8323), .ZN(n8180) );
  NAND4_X1 U7360 ( .A1(n9416), .A2(n8161), .A3(n9417), .A4(n8160), .ZN(n8162)
         );
  AND3_X1 U7361 ( .A1(n8132), .A2(n8131), .A3(n8130), .ZN(n8836) );
  NAND2_X1 U7362 ( .A1(n8165), .A2(n8164), .ZN(n7080) );
  NOR2_X1 U7363 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n7592) );
  NOR2_X1 U7364 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n7593) );
  INV_X1 U7365 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n8846) );
  INV_X4 U7366 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X4 U7367 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  XNOR2_X1 U7368 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n7480) );
  INV_X1 U7369 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n9406) );
  NOR2_X1 U7370 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n8135) );
  NOR2_X1 U7371 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n8136) );
  INV_X1 U7372 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7787) );
  NOR2_X1 U7373 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n6869) );
  NOR2_X1 U7374 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_5__SCAN_IN), .ZN(
        n6868) );
  NOR2_X1 U7375 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n6867) );
  INV_X1 U7376 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8589) );
  NOR2_X1 U7377 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n8145) );
  NOR2_X1 U7378 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n8144) );
  NAND2_X1 U7379 ( .A1(n13444), .A2(n11682), .ZN(n6424) );
  NAND2_X1 U7380 ( .A1(n13444), .A2(n11682), .ZN(n13448) );
  NOR2_X2 U7381 ( .A1(n10705), .A2(n14828), .ZN(n14737) );
  OAI22_X2 U7382 ( .A1(n10681), .A2(n10680), .B1(n10679), .B2(n6593), .ZN(
        n10928) );
  NAND2_X2 U7383 ( .A1(n10652), .A2(n10651), .ZN(n10681) );
  AOI21_X1 U7384 ( .B1(n9702), .B2(n9696), .A(n6459), .ZN(n7243) );
  NAND4_X2 U7385 ( .A1(n7635), .A2(n7634), .A3(n7633), .A4(n7632), .ZN(n12897)
         );
  NOR2_X2 U7386 ( .A1(n11695), .A2(n6648), .ZN(n11719) );
  NAND2_X1 U7387 ( .A1(n13437), .A2(n11720), .ZN(n13435) );
  INV_X4 U7388 ( .A(n9326), .ZN(n13845) );
  INV_X1 U7389 ( .A(n7545), .ZN(n7151) );
  NAND2_X1 U7390 ( .A1(n13954), .A2(n11600), .ZN(n7190) );
  INV_X1 U7391 ( .A(n12125), .ZN(n7319) );
  NOR2_X1 U7392 ( .A1(n14359), .A2(n6457), .ZN(n7247) );
  AOI21_X1 U7393 ( .B1(n6893), .B2(n6891), .A(n6495), .ZN(n6890) );
  INV_X1 U7394 ( .A(n7412), .ZN(n6891) );
  AND2_X1 U7395 ( .A1(n12889), .A2(n12890), .ZN(n12926) );
  AND2_X1 U7396 ( .A1(n7310), .A2(n7309), .ZN(n7308) );
  INV_X1 U7397 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7309) );
  INV_X1 U7398 ( .A(n7150), .ZN(n7149) );
  OAI21_X1 U7399 ( .B1(n7761), .B2(n7151), .A(n7546), .ZN(n7150) );
  AND4_X2 U7400 ( .A1(n8139), .A2(n8836), .A3(n9544), .A4(n8261), .ZN(n9592)
         );
  INV_X1 U7401 ( .A(n14578), .ZN(n11862) );
  NOR2_X1 U7402 ( .A1(n14372), .A2(n6689), .ZN(n6665) );
  INV_X1 U7403 ( .A(n7247), .ZN(n6689) );
  NOR2_X1 U7404 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n6823) );
  NOR2_X1 U7405 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n6822) );
  XNOR2_X1 U7406 ( .A(n10740), .B(SI_21_), .ZN(n10741) );
  NAND2_X1 U7407 ( .A1(n11404), .A2(n11907), .ZN(n11391) );
  NAND2_X1 U7408 ( .A1(n11455), .A2(n11442), .ZN(n12155) );
  OR2_X1 U7409 ( .A1(n14470), .A2(n11388), .ZN(n11447) );
  OR2_X1 U7410 ( .A1(n14460), .A2(n14461), .ZN(n14458) );
  AND2_X1 U7411 ( .A1(n6731), .A2(n6452), .ZN(n7503) );
  OAI21_X1 U7412 ( .B1(n12203), .B2(n12432), .A(n12202), .ZN(n12204) );
  INV_X1 U7413 ( .A(n12269), .ZN(n7397) );
  NAND2_X1 U7414 ( .A1(n7397), .A2(n6482), .ZN(n7395) );
  NAND2_X1 U7415 ( .A1(n6450), .A2(n6610), .ZN(n7145) );
  INV_X1 U7416 ( .A(n12018), .ZN(n6610) );
  INV_X1 U7417 ( .A(n12033), .ZN(n12034) );
  NAND2_X1 U7418 ( .A1(n12311), .A2(n6541), .ZN(n7385) );
  OAI21_X1 U7419 ( .B1(n13445), .B2(n12432), .A(n12322), .ZN(n12323) );
  NAND2_X1 U7420 ( .A1(n7423), .A2(n6427), .ZN(n7382) );
  INV_X1 U7421 ( .A(n7042), .ZN(n7041) );
  OAI21_X1 U7422 ( .B1(n6462), .B2(n6429), .A(n12914), .ZN(n7042) );
  OR2_X1 U7423 ( .A1(n12756), .A2(n13081), .ZN(n12918) );
  INV_X1 U7424 ( .A(n7190), .ZN(n7187) );
  AND2_X1 U7425 ( .A1(n7367), .A2(n14123), .ZN(n7366) );
  NAND2_X1 U7426 ( .A1(n7368), .A2(n11841), .ZN(n7367) );
  INV_X1 U7427 ( .A(n14204), .ZN(n7368) );
  INV_X1 U7428 ( .A(n10082), .ZN(n7331) );
  NAND2_X1 U7429 ( .A1(n8236), .A2(n8846), .ZN(n6605) );
  NAND2_X1 U7430 ( .A1(n6579), .A2(n7431), .ZN(n7432) );
  NAND2_X1 U7431 ( .A1(n7477), .A2(n7430), .ZN(n6579) );
  INV_X1 U7432 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7430) );
  INV_X1 U7433 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7591) );
  INV_X1 U7434 ( .A(n6885), .ZN(n6884) );
  AOI21_X1 U7435 ( .B1(n7015), .B2(n7017), .A(n7014), .ZN(n7013) );
  INV_X1 U7436 ( .A(n12880), .ZN(n7014) );
  OR2_X1 U7437 ( .A1(n12535), .A2(n12538), .ZN(n12858) );
  AND2_X1 U7438 ( .A1(n12830), .A2(n12831), .ZN(n12938) );
  INV_X1 U7439 ( .A(n10042), .ZN(n12773) );
  OAI21_X1 U7440 ( .B1(n8099), .B2(n8098), .A(n8899), .ZN(n8120) );
  INV_X1 U7441 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8104) );
  INV_X1 U7442 ( .A(n7789), .ZN(n6704) );
  NOR2_X1 U7443 ( .A1(n13964), .A2(n13973), .ZN(n6954) );
  NAND2_X1 U7444 ( .A1(n6966), .A2(n6965), .ZN(n13597) );
  AOI21_X1 U7445 ( .B1(n6968), .B2(n6970), .A(n6477), .ZN(n6965) );
  INV_X1 U7446 ( .A(n7192), .ZN(n7185) );
  AND2_X1 U7447 ( .A1(n9486), .A2(n9481), .ZN(n6979) );
  AOI21_X1 U7448 ( .B1(n6930), .B2(n6934), .A(n6928), .ZN(n6927) );
  NAND2_X1 U7449 ( .A1(n10186), .A2(n6930), .ZN(n6929) );
  NOR2_X1 U7450 ( .A1(n10740), .A2(SI_21_), .ZN(n6928) );
  OR2_X1 U7451 ( .A1(n8380), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8629) );
  INV_X1 U7452 ( .A(n6558), .ZN(n6852) );
  INV_X1 U7453 ( .A(n11935), .ZN(n8704) );
  INV_X1 U7454 ( .A(n8693), .ZN(n8695) );
  NOR2_X1 U7455 ( .A1(n12103), .A2(n14566), .ZN(n6805) );
  NAND2_X1 U7456 ( .A1(n7069), .A2(n6464), .ZN(n7068) );
  NAND2_X1 U7457 ( .A1(n7070), .A2(n7072), .ZN(n7069) );
  NOR2_X1 U7458 ( .A1(n14430), .A2(n6777), .ZN(n6776) );
  INV_X1 U7459 ( .A(n6779), .ZN(n6777) );
  NAND2_X1 U7460 ( .A1(n12039), .A2(n6433), .ZN(n6785) );
  NOR2_X1 U7461 ( .A1(n11356), .A2(n7267), .ZN(n7266) );
  INV_X1 U7462 ( .A(n11352), .ZN(n7267) );
  AND2_X1 U7463 ( .A1(n14514), .A2(n11443), .ZN(n7096) );
  NOR2_X1 U7464 ( .A1(n10548), .A2(n7261), .ZN(n7260) );
  INV_X1 U7465 ( .A(n10547), .ZN(n7261) );
  NAND2_X1 U7466 ( .A1(n8710), .A2(n12110), .ZN(n11935) );
  NAND2_X1 U7467 ( .A1(n7245), .A2(n14344), .ZN(n6664) );
  INV_X1 U7468 ( .A(n11931), .ZN(n8710) );
  NOR2_X1 U7469 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n9419) );
  AOI21_X1 U7470 ( .B1(n11330), .B2(n7339), .A(n7336), .ZN(n7335) );
  INV_X1 U7471 ( .A(n11291), .ZN(n7336) );
  INV_X1 U7472 ( .A(n6600), .ZN(n6599) );
  OAI21_X1 U7473 ( .B1(n11158), .B2(n6924), .A(n6916), .ZN(n6600) );
  OAI21_X1 U7474 ( .B1(n11158), .B2(n6922), .A(n6920), .ZN(n6918) );
  INV_X1 U7475 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U7476 ( .A1(n6571), .A2(n9540), .ZN(n9584) );
  XNOR2_X1 U7477 ( .A(n7432), .B(n6820), .ZN(n7476) );
  INV_X1 U7478 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n6820) );
  OAI21_X1 U7479 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n7445), .A(n7444), .ZN(
        n7474) );
  XNOR2_X1 U7480 ( .A(n7165), .B(n9776), .ZN(n12953) );
  INV_X1 U7481 ( .A(n7404), .ZN(n7168) );
  INV_X1 U7482 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7590) );
  XNOR2_X1 U7483 ( .A(n11115), .B(n11121), .ZN(n10793) );
  AND2_X1 U7484 ( .A1(n12914), .A2(n11654), .ZN(n12949) );
  NOR2_X1 U7485 ( .A1(n12947), .A2(n6717), .ZN(n6716) );
  INV_X1 U7486 ( .A(n8026), .ZN(n6717) );
  AND2_X1 U7487 ( .A1(n12763), .A2(n7992), .ZN(n13148) );
  NAND2_X1 U7488 ( .A1(n13232), .A2(n6904), .ZN(n6900) );
  AOI21_X1 U7489 ( .B1(n7034), .B2(n7032), .A(n7031), .ZN(n7030) );
  INV_X1 U7490 ( .A(n12852), .ZN(n7031) );
  NOR2_X1 U7491 ( .A1(n6453), .A2(n13249), .ZN(n7032) );
  NAND2_X1 U7492 ( .A1(n7034), .A2(n12942), .ZN(n7033) );
  OR2_X1 U7493 ( .A1(n8119), .A2(n12761), .ZN(n14762) );
  INV_X1 U7494 ( .A(n7749), .ZN(n12748) );
  NAND2_X1 U7495 ( .A1(n7173), .A2(n7174), .ZN(n12503) );
  AOI21_X1 U7496 ( .B1(n7175), .B2(n11648), .A(n6559), .ZN(n7174) );
  AND2_X1 U7497 ( .A1(n7606), .A2(n7595), .ZN(n7058) );
  NOR2_X2 U7498 ( .A1(n7603), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n7614) );
  NAND2_X1 U7499 ( .A1(n7584), .A2(n11163), .ZN(n7172) );
  CLKBUF_X1 U7500 ( .A(n8968), .Z(n6772) );
  NAND2_X1 U7501 ( .A1(n7959), .A2(n7576), .ZN(n7969) );
  AOI21_X1 U7502 ( .B1(n7940), .B2(n7158), .A(n7157), .ZN(n7156) );
  INV_X1 U7503 ( .A(n7570), .ZN(n7157) );
  INV_X1 U7504 ( .A(n7568), .ZN(n7158) );
  INV_X1 U7505 ( .A(n7940), .ZN(n7159) );
  INV_X1 U7506 ( .A(n7895), .ZN(n7164) );
  XNOR2_X1 U7507 ( .A(n12281), .B(n6627), .ZN(n10406) );
  XNOR2_X1 U7508 ( .A(n12245), .B(n13459), .ZN(n9703) );
  XNOR2_X1 U7509 ( .A(n9602), .B(n7226), .ZN(n7228) );
  INV_X1 U7510 ( .A(n9106), .ZN(n7226) );
  XNOR2_X1 U7511 ( .A(n13459), .B(n12194), .ZN(n9602) );
  NAND2_X1 U7512 ( .A1(n10719), .A2(n10718), .ZN(n11067) );
  AND2_X1 U7513 ( .A1(n14076), .A2(n14073), .ZN(n8853) );
  AND2_X1 U7514 ( .A1(n8593), .A2(n6960), .ZN(n11528) );
  AND2_X1 U7515 ( .A1(n11588), .A2(n11589), .ZN(n13791) );
  NAND2_X1 U7516 ( .A1(n10700), .A2(n10699), .ZN(n10921) );
  OAI21_X1 U7517 ( .B1(n10567), .B2(n6987), .A(n6988), .ZN(n10700) );
  AND2_X1 U7518 ( .A1(n6990), .A2(n6989), .ZN(n6988) );
  NAND2_X1 U7519 ( .A1(n10567), .A2(n10566), .ZN(n6993) );
  NAND2_X1 U7520 ( .A1(n12460), .A2(n7196), .ZN(n7195) );
  INV_X1 U7521 ( .A(n9764), .ZN(n7196) );
  NAND2_X1 U7522 ( .A1(n9909), .A2(n9908), .ZN(n10238) );
  NAND2_X1 U7523 ( .A1(n8931), .A2(n11907), .ZN(n8848) );
  NAND2_X1 U7524 ( .A1(n8931), .A2(n8968), .ZN(n8843) );
  CLKBUF_X1 U7525 ( .A(n8602), .Z(n13603) );
  INV_X1 U7526 ( .A(n13947), .ZN(n6660) );
  CLKBUF_X3 U7527 ( .A(n8848), .Z(n12399) );
  NAND2_X1 U7528 ( .A1(n9592), .A2(n6662), .ZN(n8585) );
  AND2_X1 U7529 ( .A1(n6420), .A2(n6518), .ZN(n6662) );
  AND2_X1 U7530 ( .A1(n6420), .A2(n7214), .ZN(n7212) );
  NOR2_X1 U7531 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n7214) );
  INV_X1 U7532 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8138) );
  OR2_X1 U7533 ( .A1(n6853), .A2(n6852), .ZN(n6850) );
  AND2_X1 U7534 ( .A1(n9614), .A2(n10109), .ZN(n6853) );
  OR2_X1 U7535 ( .A1(n6852), .A2(n7406), .ZN(n6851) );
  AOI21_X1 U7536 ( .B1(n7362), .B2(n7364), .A(n6507), .ZN(n7360) );
  AOI21_X1 U7537 ( .B1(n7360), .B2(n6843), .A(n6539), .ZN(n6842) );
  INV_X1 U7538 ( .A(n7362), .ZN(n6843) );
  AND2_X1 U7539 ( .A1(n11917), .A2(n11935), .ZN(n11793) );
  NOR2_X1 U7540 ( .A1(n7109), .A2(n7107), .ZN(n7106) );
  INV_X1 U7541 ( .A(n12173), .ZN(n7109) );
  NAND2_X2 U7542 ( .A1(n8696), .A2(n8695), .ZN(n11435) );
  INV_X1 U7543 ( .A(n8996), .ZN(n11921) );
  AOI21_X1 U7544 ( .B1(n11446), .B2(n12044), .A(n7410), .ZN(n14457) );
  AND2_X1 U7545 ( .A1(n11447), .A2(n11389), .ZN(n14461) );
  AND2_X1 U7546 ( .A1(n12140), .A2(n10525), .ZN(n7093) );
  OR2_X1 U7547 ( .A1(n8784), .A2(n8710), .ZN(n8807) );
  AND3_X1 U7548 ( .A1(n8344), .A2(n8347), .A3(n8343), .ZN(n8780) );
  OR2_X1 U7549 ( .A1(n12113), .A2(n12112), .ZN(n12115) );
  AND3_X1 U7550 ( .A1(n6825), .A2(n6824), .A3(n8180), .ZN(n7078) );
  INV_X1 U7551 ( .A(n7080), .ZN(n6825) );
  AND2_X1 U7552 ( .A1(n8336), .A2(n8179), .ZN(n6824) );
  OAI21_X1 U7553 ( .B1(n8834), .B2(n6940), .A(n6938), .ZN(n9537) );
  NAND2_X1 U7554 ( .A1(n7450), .A2(n7449), .ZN(n7472) );
  OR2_X1 U7555 ( .A1(n7509), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n7449) );
  NOR2_X2 U7556 ( .A1(n15193), .A2(n12771), .ZN(n15190) );
  AND2_X1 U7557 ( .A1(n9120), .A2(n9112), .ZN(n7232) );
  NAND2_X1 U7558 ( .A1(n11393), .A2(n11392), .ZN(n14451) );
  NAND2_X1 U7559 ( .A1(n14824), .A2(n7372), .ZN(n11208) );
  NOR2_X1 U7560 ( .A1(n11032), .A2(n7373), .ZN(n7372) );
  INV_X1 U7561 ( .A(n11026), .ZN(n7373) );
  XNOR2_X1 U7562 ( .A(n6621), .B(n6620), .ZN(n14565) );
  INV_X1 U7563 ( .A(n12157), .ZN(n6620) );
  NAND2_X1 U7564 ( .A1(n14566), .A2(n14345), .ZN(n6622) );
  INV_X1 U7565 ( .A(n7504), .ZN(n6808) );
  INV_X1 U7566 ( .A(n7521), .ZN(n6809) );
  OAI21_X1 U7567 ( .B1(n12197), .B2(n12196), .A(n12195), .ZN(n12199) );
  NAND2_X1 U7568 ( .A1(n6695), .A2(n6698), .ZN(n12222) );
  INV_X1 U7569 ( .A(n12216), .ZN(n6677) );
  OR2_X1 U7570 ( .A1(n7124), .A2(n11978), .ZN(n7126) );
  AOI21_X1 U7571 ( .B1(n11978), .B2(n7124), .A(n7125), .ZN(n7123) );
  INV_X1 U7572 ( .A(n11986), .ZN(n7131) );
  NAND2_X1 U7573 ( .A1(n7390), .A2(n6443), .ZN(n7389) );
  INV_X1 U7574 ( .A(n12250), .ZN(n6685) );
  AOI21_X1 U7575 ( .B1(n7396), .B2(n7395), .A(n6520), .ZN(n7394) );
  NOR2_X1 U7576 ( .A1(n7397), .A2(n6482), .ZN(n7396) );
  NAND2_X1 U7577 ( .A1(n7145), .A2(n12028), .ZN(n7143) );
  INV_X1 U7578 ( .A(n12282), .ZN(n6675) );
  INV_X1 U7579 ( .A(n12283), .ZN(n6616) );
  INV_X1 U7580 ( .A(n12284), .ZN(n6617) );
  INV_X1 U7581 ( .A(n12043), .ZN(n7141) );
  NAND2_X1 U7582 ( .A1(n6567), .A2(n6566), .ZN(n6631) );
  INV_X1 U7583 ( .A(n12296), .ZN(n6566) );
  AOI22_X1 U7584 ( .A1(n12314), .A2(n12408), .B1(n13545), .B2(n12403), .ZN(
        n12315) );
  INV_X1 U7585 ( .A(n12065), .ZN(n7132) );
  NOR2_X1 U7586 ( .A1(n7134), .A2(n12065), .ZN(n7133) );
  NAND2_X1 U7587 ( .A1(n7392), .A2(n6481), .ZN(n7391) );
  NAND2_X1 U7588 ( .A1(n6548), .A2(n12344), .ZN(n7400) );
  NAND2_X1 U7589 ( .A1(n11916), .A2(n11917), .ZN(n7112) );
  INV_X1 U7590 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7599) );
  INV_X1 U7591 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7656) );
  NAND2_X1 U7592 ( .A1(n6572), .A2(n6487), .ZN(n7379) );
  INV_X1 U7593 ( .A(n12354), .ZN(n6572) );
  INV_X1 U7594 ( .A(n12353), .ZN(n7380) );
  NAND2_X1 U7595 ( .A1(n6517), .A2(n7382), .ZN(n7381) );
  AND2_X1 U7596 ( .A1(n11473), .A2(n12488), .ZN(n12181) );
  NOR2_X1 U7597 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n8132) );
  NOR2_X1 U7598 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8130) );
  NOR2_X1 U7599 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8131) );
  NOR2_X1 U7600 ( .A1(n7089), .A2(n9939), .ZN(n7088) );
  INV_X1 U7601 ( .A(n9684), .ZN(n7089) );
  NOR2_X1 U7602 ( .A1(n11289), .A2(SI_25_), .ZN(n7340) );
  INV_X1 U7603 ( .A(n11159), .ZN(n6922) );
  INV_X1 U7604 ( .A(n6921), .ZN(n6920) );
  OAI21_X1 U7605 ( .B1(n11157), .B2(n6922), .A(SI_24_), .ZN(n6921) );
  INV_X1 U7606 ( .A(n7330), .ZN(n7329) );
  OAI21_X1 U7607 ( .B1(n10077), .B2(n7331), .A(n10179), .ZN(n7330) );
  AOI21_X1 U7608 ( .B1(n6938), .B2(n6940), .A(n6937), .ZN(n6936) );
  INV_X1 U7609 ( .A(n9536), .ZN(n6937) );
  INV_X1 U7610 ( .A(n9409), .ZN(n9414) );
  INV_X1 U7611 ( .A(n7347), .ZN(n7346) );
  AND2_X1 U7612 ( .A1(n7348), .A2(n9031), .ZN(n7347) );
  INV_X1 U7613 ( .A(n9036), .ZN(n7348) );
  INV_X1 U7614 ( .A(n13222), .ZN(n12538) );
  INV_X1 U7615 ( .A(n12543), .ZN(n7299) );
  AOI21_X1 U7616 ( .B1(n11655), .B2(n7041), .A(n7038), .ZN(n7037) );
  NAND2_X1 U7617 ( .A1(n7039), .A2(n12754), .ZN(n7038) );
  NAND2_X1 U7618 ( .A1(n7041), .A2(n6429), .ZN(n7039) );
  OR2_X1 U7619 ( .A1(n12564), .A2(n12565), .ZN(n12893) );
  AND2_X1 U7620 ( .A1(n12766), .A2(n12890), .ZN(n7055) );
  OR2_X1 U7621 ( .A1(n12695), .A2(n13175), .ZN(n12880) );
  INV_X1 U7622 ( .A(n6904), .ZN(n6898) );
  NOR2_X1 U7623 ( .A1(n13225), .A2(n13237), .ZN(n6904) );
  AND2_X1 U7624 ( .A1(n6901), .A2(n13214), .ZN(n6899) );
  INV_X1 U7625 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7606) );
  INV_X1 U7626 ( .A(n7578), .ZN(n7182) );
  INV_X1 U7627 ( .A(n7968), .ZN(n7179) );
  NOR2_X1 U7628 ( .A1(n7929), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n7659) );
  AOI21_X1 U7629 ( .B1(n13448), .B2(n6765), .A(n6761), .ZN(n11693) );
  INV_X1 U7630 ( .A(n13830), .ZN(n11627) );
  AND2_X1 U7631 ( .A1(n13820), .A2(n6984), .ZN(n6983) );
  NAND2_X1 U7632 ( .A1(n13841), .A2(n11639), .ZN(n6984) );
  INV_X1 U7633 ( .A(n13803), .ZN(n7202) );
  INV_X1 U7634 ( .A(n11549), .ZN(n7203) );
  INV_X1 U7635 ( .A(n10568), .ZN(n6992) );
  NOR2_X1 U7636 ( .A1(n9761), .A2(n12259), .ZN(n6951) );
  OR2_X1 U7637 ( .A1(n14006), .A2(n11242), .ZN(n13898) );
  OAI21_X1 U7638 ( .B1(n8141), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8153) );
  NAND2_X1 U7639 ( .A1(n14068), .A2(n6657), .ZN(n6656) );
  NAND2_X1 U7640 ( .A1(n8573), .A2(n6657), .ZN(n8491) );
  NOR2_X1 U7641 ( .A1(n11449), .A2(n7252), .ZN(n7251) );
  INV_X1 U7642 ( .A(n7256), .ZN(n7252) );
  NOR2_X1 U7643 ( .A1(n12149), .A2(n6788), .ZN(n6787) );
  INV_X1 U7644 ( .A(n12024), .ZN(n6788) );
  AND2_X1 U7645 ( .A1(n12133), .A2(n7090), .ZN(n7086) );
  NAND2_X1 U7646 ( .A1(n14262), .A2(n7091), .ZN(n7090) );
  NAND2_X1 U7647 ( .A1(n9685), .A2(n7088), .ZN(n7087) );
  OR2_X1 U7648 ( .A1(n14264), .A2(n14938), .ZN(n11957) );
  NAND2_X1 U7649 ( .A1(n7343), .A2(n7342), .ZN(n7341) );
  INV_X1 U7650 ( .A(n7340), .ZN(n7338) );
  NAND2_X1 U7651 ( .A1(n9028), .A2(n9027), .ZN(n7349) );
  NAND2_X1 U7652 ( .A1(n7349), .A2(n7347), .ZN(n9412) );
  NAND4_X1 U7653 ( .A1(n13069), .A2(n7312), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7311) );
  INV_X1 U7654 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7315) );
  AND2_X1 U7655 ( .A1(n7483), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n7481) );
  NAND2_X1 U7656 ( .A1(n6815), .A2(n6813), .ZN(n7429) );
  NAND2_X1 U7657 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n6814), .ZN(n6813) );
  INV_X1 U7658 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6814) );
  XNOR2_X1 U7659 ( .A(n7434), .B(n6818), .ZN(n7489) );
  INV_X1 U7660 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n6818) );
  NOR2_X1 U7661 ( .A1(n10056), .A2(n15194), .ZN(n7275) );
  NOR2_X1 U7662 ( .A1(n10060), .A2(n7275), .ZN(n7274) );
  NAND2_X1 U7663 ( .A1(n7278), .A2(n7277), .ZN(n7276) );
  INV_X1 U7664 ( .A(n10058), .ZN(n7278) );
  NAND2_X1 U7665 ( .A1(n7288), .A2(n7287), .ZN(n12613) );
  AOI21_X1 U7666 ( .B1(n7290), .B2(n7292), .A(n6542), .ZN(n7287) );
  NAND2_X1 U7667 ( .A1(n12640), .A2(n7290), .ZN(n7288) );
  NAND2_X1 U7668 ( .A1(n6888), .A2(n7702), .ZN(n9779) );
  INV_X1 U7669 ( .A(n6889), .ZN(n6888) );
  NAND2_X1 U7670 ( .A1(n8005), .A2(SI_1_), .ZN(n7702) );
  NOR2_X1 U7671 ( .A1(n12623), .A2(n7302), .ZN(n7301) );
  INV_X1 U7672 ( .A(n12546), .ZN(n7302) );
  AOI21_X1 U7673 ( .B1(n12691), .B2(n13175), .A(n12552), .ZN(n12555) );
  NOR2_X1 U7674 ( .A1(n12549), .A2(n12551), .ZN(n12552) );
  INV_X1 U7675 ( .A(n7274), .ZN(n7270) );
  NAND2_X1 U7676 ( .A1(n10089), .A2(n15172), .ZN(n7279) );
  NAND2_X1 U7677 ( .A1(n12709), .A2(n12536), .ZN(n12672) );
  INV_X1 U7678 ( .A(n12594), .ZN(n7307) );
  INV_X1 U7679 ( .A(n12522), .ZN(n7306) );
  INV_X1 U7680 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8030) );
  INV_X1 U7681 ( .A(n7730), .ZN(n7296) );
  NAND2_X1 U7682 ( .A1(n7591), .A2(n6866), .ZN(n7297) );
  INV_X1 U7683 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n6866) );
  NAND2_X1 U7684 ( .A1(n6755), .A2(n6753), .ZN(n10158) );
  NAND2_X1 U7685 ( .A1(n15115), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n6755) );
  NAND2_X1 U7686 ( .A1(n6754), .A2(n15127), .ZN(n6753) );
  NAND2_X1 U7687 ( .A1(n9962), .A2(n9963), .ZN(n6754) );
  NAND2_X1 U7688 ( .A1(n6758), .A2(n6757), .ZN(n10336) );
  NAND2_X1 U7689 ( .A1(n15135), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n6757) );
  OAI21_X1 U7690 ( .B1(n15135), .B2(P3_REG2_REG_8__SCAN_IN), .A(n15149), .ZN(
        n6758) );
  NAND2_X1 U7691 ( .A1(n12988), .A2(n10792), .ZN(n11115) );
  NAND2_X1 U7692 ( .A1(n10793), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n11116) );
  XNOR2_X1 U7693 ( .A(n12899), .B(n12897), .ZN(n12947) );
  INV_X1 U7694 ( .A(n8002), .ZN(n6724) );
  NAND2_X1 U7695 ( .A1(n13134), .A2(n7412), .ZN(n6894) );
  AND2_X1 U7696 ( .A1(n12880), .A2(n6471), .ZN(n13165) );
  NAND2_X1 U7697 ( .A1(n6431), .A2(n12873), .ZN(n7018) );
  NAND2_X1 U7698 ( .A1(n7019), .A2(n6431), .ZN(n7017) );
  NAND2_X1 U7699 ( .A1(n13189), .A2(n13188), .ZN(n13187) );
  OAI21_X1 U7700 ( .B1(n13226), .B2(n7046), .A(n7044), .ZN(n7049) );
  AOI21_X1 U7701 ( .B1(n7045), .B2(n7047), .A(n8059), .ZN(n7044) );
  INV_X1 U7702 ( .A(n7047), .ZN(n7046) );
  AND2_X1 U7703 ( .A1(n6903), .A2(n6902), .ZN(n6901) );
  OR2_X1 U7704 ( .A1(n13322), .A2(n13234), .ZN(n6902) );
  OR2_X1 U7705 ( .A1(n13225), .A2(n6906), .ZN(n6903) );
  NOR2_X1 U7706 ( .A1(n13214), .A2(n7048), .ZN(n7047) );
  NAND2_X1 U7707 ( .A1(n13226), .A2(n13225), .ZN(n13224) );
  AND2_X1 U7708 ( .A1(n12857), .A2(n12860), .ZN(n13225) );
  OR2_X1 U7709 ( .A1(n13380), .A2(n13235), .ZN(n7413) );
  AOI21_X1 U7710 ( .B1(n7030), .B2(n7033), .A(n13231), .ZN(n7027) );
  AND2_X1 U7711 ( .A1(n6876), .A2(n6440), .ZN(n6874) );
  AND2_X1 U7712 ( .A1(n13260), .A2(n6877), .ZN(n6876) );
  NAND2_X1 U7713 ( .A1(n14755), .A2(n6878), .ZN(n6877) );
  NAND2_X1 U7714 ( .A1(n6516), .A2(n12843), .ZN(n7034) );
  AND2_X1 U7715 ( .A1(n12844), .A2(n12843), .ZN(n13266) );
  AOI21_X1 U7716 ( .B1(n7052), .B2(n10886), .A(n7051), .ZN(n7050) );
  INV_X1 U7717 ( .A(n12827), .ZN(n7051) );
  INV_X1 U7718 ( .A(n15192), .ZN(n14778) );
  NAND2_X1 U7719 ( .A1(n8055), .A2(n12927), .ZN(n10880) );
  NAND2_X1 U7720 ( .A1(n10817), .A2(n6909), .ZN(n10884) );
  NOR2_X1 U7721 ( .A1(n6911), .A2(n6910), .ZN(n6909) );
  INV_X1 U7722 ( .A(n7889), .ZN(n6910) );
  INV_X1 U7723 ( .A(n7890), .ZN(n6911) );
  AND2_X1 U7724 ( .A1(n10817), .A2(n7889), .ZN(n10881) );
  INV_X1 U7725 ( .A(n12932), .ZN(n10812) );
  AND2_X1 U7726 ( .A1(n8046), .A2(n12917), .ZN(n15195) );
  NAND2_X1 U7727 ( .A1(n9799), .A2(n9798), .ZN(n9802) );
  NAND2_X1 U7728 ( .A1(n13394), .A2(n12748), .ZN(n12747) );
  OR2_X1 U7729 ( .A1(n13081), .A2(n13080), .ZN(n13335) );
  INV_X1 U7730 ( .A(n11898), .ZN(n6709) );
  NAND2_X1 U7731 ( .A1(n11659), .A2(n11658), .ZN(n13277) );
  INV_X1 U7732 ( .A(n14762), .ZN(n15198) );
  INV_X1 U7733 ( .A(n15195), .ZN(n14776) );
  NAND2_X1 U7734 ( .A1(n12962), .A2(n10042), .ZN(n15226) );
  INV_X1 U7735 ( .A(n8087), .ZN(n8899) );
  OAI21_X1 U7736 ( .B1(n8015), .B2(n7587), .A(n7588), .ZN(n11649) );
  XNOR2_X1 U7737 ( .A(n8078), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8086) );
  NOR2_X1 U7738 ( .A1(n11565), .A2(n6722), .ZN(n6721) );
  INV_X1 U7739 ( .A(n7579), .ZN(n6722) );
  MUX2_X1 U7740 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8072), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8073) );
  NAND2_X1 U7741 ( .A1(n7969), .A2(n7968), .ZN(n7971) );
  NAND2_X1 U7742 ( .A1(n7575), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7576) );
  NAND2_X1 U7743 ( .A1(n7659), .A2(n7945), .ZN(n7668) );
  AND2_X1 U7744 ( .A1(n7572), .A2(n7571), .ZN(n7664) );
  NAND2_X1 U7745 ( .A1(n7155), .A2(n7153), .ZN(n7667) );
  AOI21_X1 U7746 ( .B1(n7156), .B2(n7159), .A(n7154), .ZN(n7153) );
  NAND2_X1 U7747 ( .A1(n7928), .A2(n7156), .ZN(n7155) );
  INV_X1 U7748 ( .A(n7664), .ZN(n7154) );
  INV_X1 U7749 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7945) );
  AND2_X1 U7750 ( .A1(n7570), .A2(n7569), .ZN(n7940) );
  NAND2_X1 U7751 ( .A1(n7912), .A2(n7566), .ZN(n7926) );
  AND2_X1 U7752 ( .A1(n7568), .A2(n7567), .ZN(n7925) );
  NAND2_X1 U7753 ( .A1(n7926), .A2(n7925), .ZN(n7928) );
  OAI21_X1 U7754 ( .B1(n7562), .B2(n7164), .A(n7564), .ZN(n7163) );
  NAND2_X1 U7755 ( .A1(n6711), .A2(n7160), .ZN(n7912) );
  NAND2_X1 U7756 ( .A1(n7680), .A2(n7162), .ZN(n6711) );
  AOI21_X1 U7757 ( .B1(n7162), .B2(n7164), .A(n7161), .ZN(n7160) );
  INV_X1 U7758 ( .A(n7909), .ZN(n7161) );
  AND2_X1 U7759 ( .A1(n7564), .A2(n7563), .ZN(n7895) );
  OR2_X1 U7760 ( .A1(n7560), .A2(n9039), .ZN(n7561) );
  NAND2_X1 U7761 ( .A1(n7560), .A2(n9039), .ZN(n7562) );
  NAND2_X1 U7762 ( .A1(n6712), .A2(n7561), .ZN(n7680) );
  AND2_X1 U7763 ( .A1(n7562), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n6712) );
  INV_X1 U7764 ( .A(n6702), .ZN(n6701) );
  OAI21_X1 U7765 ( .B1(n6455), .B2(n6703), .A(n7811), .ZN(n6702) );
  INV_X1 U7766 ( .A(n7548), .ZN(n6703) );
  AOI21_X1 U7767 ( .B1(n7149), .B2(n7151), .A(n6509), .ZN(n7147) );
  NAND2_X1 U7768 ( .A1(n7762), .A2(n7149), .ZN(n7146) );
  NAND2_X1 U7769 ( .A1(n7146), .A2(n6455), .ZN(n7792) );
  AND2_X1 U7770 ( .A1(n7545), .A2(n7544), .ZN(n7761) );
  NAND2_X1 U7771 ( .A1(n6700), .A2(n7540), .ZN(n7748) );
  XNOR2_X1 U7772 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7534) );
  NAND2_X1 U7773 ( .A1(n10653), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n10686) );
  INV_X1 U7774 ( .A(n10654), .ZN(n10653) );
  OR2_X1 U7775 ( .A1(n10934), .A2(n11084), .ZN(n11075) );
  XNOR2_X1 U7776 ( .A(n12259), .B(n13459), .ZN(n9844) );
  NAND2_X1 U7777 ( .A1(n10410), .A2(n10409), .ZN(n10416) );
  XNOR2_X1 U7778 ( .A(n12268), .B(n6627), .ZN(n11742) );
  NAND2_X1 U7779 ( .A1(n7237), .A2(n11734), .ZN(n7236) );
  INV_X1 U7780 ( .A(n7239), .ZN(n7237) );
  NOR2_X1 U7781 ( .A1(n7239), .A2(n11733), .ZN(n7238) );
  INV_X1 U7782 ( .A(n8853), .ZN(n8942) );
  AND2_X1 U7783 ( .A1(n8595), .A2(n8596), .ZN(n6615) );
  NAND2_X1 U7784 ( .A1(n6591), .A2(n8507), .ZN(n8618) );
  OR2_X1 U7785 ( .A1(n15047), .A2(n15048), .ZN(n6641) );
  NOR2_X1 U7786 ( .A1(n10457), .A2(n6642), .ZN(n10624) );
  AND2_X1 U7787 ( .A1(n10648), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6642) );
  AND2_X1 U7788 ( .A1(n12479), .A2(n11643), .ZN(n6972) );
  NAND2_X1 U7789 ( .A1(n12479), .A2(n6504), .ZN(n6971) );
  INV_X1 U7790 ( .A(n12478), .ZN(n6973) );
  NAND2_X1 U7791 ( .A1(n13780), .A2(n13536), .ZN(n7192) );
  NAND2_X1 U7792 ( .A1(n11641), .A2(n11640), .ZN(n13792) );
  AND2_X1 U7793 ( .A1(n11563), .A2(n13803), .ZN(n13827) );
  NAND2_X1 U7794 ( .A1(n6986), .A2(n6985), .ZN(n13838) );
  INV_X1 U7795 ( .A(n13841), .ZN(n6985) );
  AND2_X1 U7796 ( .A1(n11535), .A2(n11524), .ZN(n7218) );
  AND2_X1 U7797 ( .A1(n11502), .A2(n11501), .ZN(n13890) );
  INV_X1 U7798 ( .A(n13896), .ZN(n6999) );
  NAND2_X1 U7799 ( .A1(n11224), .A2(n11223), .ZN(n11634) );
  NAND2_X1 U7800 ( .A1(n10931), .A2(n6493), .ZN(n11142) );
  AND2_X1 U7801 ( .A1(n12471), .A2(n10922), .ZN(n7003) );
  OR2_X1 U7802 ( .A1(n10921), .A2(n10920), .ZN(n7004) );
  OR2_X1 U7803 ( .A1(n14017), .A2(n13549), .ZN(n6994) );
  NAND2_X1 U7804 ( .A1(n10359), .A2(n7222), .ZN(n10559) );
  AND2_X1 U7805 ( .A1(n12466), .A2(n10358), .ZN(n7222) );
  NAND2_X1 U7806 ( .A1(n10371), .A2(n10370), .ZN(n10567) );
  NAND2_X1 U7807 ( .A1(n6951), .A2(n6950), .ZN(n10252) );
  AOI21_X1 U7808 ( .B1(n6430), .B2(n7197), .A(n10237), .ZN(n7193) );
  OAI21_X1 U7809 ( .B1(n9435), .B2(n6978), .A(n6976), .ZN(n9907) );
  AOI21_X1 U7810 ( .B1(n6979), .B2(n6977), .A(n6480), .ZN(n6976) );
  INV_X1 U7811 ( .A(n6979), .ZN(n6978) );
  NAND2_X1 U7812 ( .A1(n7207), .A2(n6437), .ZN(n9487) );
  NAND2_X1 U7813 ( .A1(n9435), .A2(n12458), .ZN(n9482) );
  NAND2_X1 U7814 ( .A1(n10312), .A2(n12456), .ZN(n10311) );
  XNOR2_X1 U7815 ( .A(n12194), .B(n13561), .ZN(n8680) );
  OR2_X1 U7816 ( .A1(n9089), .A2(n9092), .ZN(n9124) );
  NAND2_X1 U7817 ( .A1(n12396), .A2(n12395), .ZN(n13579) );
  NAND2_X1 U7818 ( .A1(n11605), .A2(n11604), .ZN(n13944) );
  AND2_X1 U7819 ( .A1(n13599), .A2(n13598), .ZN(n13949) );
  OR2_X1 U7820 ( .A1(n13597), .A2(n13596), .ZN(n13598) );
  OAI21_X1 U7821 ( .B1(n13772), .B2(n7189), .A(n7183), .ZN(n13592) );
  NOR2_X1 U7822 ( .A1(n6434), .A2(n6425), .ZN(n7183) );
  NAND2_X1 U7823 ( .A1(n11492), .A2(n11491), .ZN(n13960) );
  AND2_X1 U7824 ( .A1(n10826), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8578) );
  NOR2_X1 U7825 ( .A1(n8585), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n6964) );
  AND2_X1 U7826 ( .A1(n6420), .A2(n13732), .ZN(n7213) );
  INV_X1 U7827 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n13732) );
  NAND2_X1 U7828 ( .A1(n10745), .A2(n7352), .ZN(n7351) );
  OR2_X1 U7829 ( .A1(n10744), .A2(n10743), .ZN(n10798) );
  INV_X1 U7830 ( .A(n9593), .ZN(n10075) );
  AND2_X1 U7831 ( .A1(n8381), .A2(n8629), .ZN(n9705) );
  AND2_X1 U7832 ( .A1(n8262), .A2(n8261), .ZN(n8837) );
  INV_X1 U7833 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8598) );
  OR2_X1 U7834 ( .A1(n14177), .A2(n6831), .ZN(n6830) );
  AOI21_X1 U7835 ( .B1(n6842), .B2(n6844), .A(n6497), .ZN(n6840) );
  INV_X1 U7836 ( .A(n7360), .ZN(n6844) );
  AOI21_X1 U7837 ( .B1(n6850), .B2(n6851), .A(n6848), .ZN(n6847) );
  INV_X1 U7838 ( .A(n14093), .ZN(n6848) );
  INV_X1 U7839 ( .A(n14254), .ZN(n11212) );
  NAND3_X1 U7840 ( .A1(n14230), .A2(n11799), .A3(n11795), .ZN(n14165) );
  AOI21_X1 U7841 ( .B1(n6861), .B2(n6863), .A(n6859), .ZN(n6858) );
  INV_X1 U7842 ( .A(n7365), .ZN(n6859) );
  NOR2_X1 U7843 ( .A1(n10979), .A2(n10978), .ZN(n11172) );
  OR2_X1 U7844 ( .A1(n11919), .A2(n8788), .ZN(n8790) );
  AND2_X1 U7845 ( .A1(n8791), .A2(n8789), .ZN(n6561) );
  NAND2_X1 U7846 ( .A1(n11915), .A2(n11914), .ZN(n12159) );
  NAND2_X1 U7847 ( .A1(n12118), .A2(n12117), .ZN(n14331) );
  NAND2_X1 U7848 ( .A1(n6601), .A2(n11913), .ZN(n12118) );
  INV_X1 U7849 ( .A(n14074), .ZN(n6601) );
  NAND2_X1 U7850 ( .A1(n11300), .A2(n11299), .ZN(n12103) );
  OAI21_X1 U7851 ( .B1(n14360), .B2(n7068), .A(n7066), .ZN(n11758) );
  INV_X1 U7852 ( .A(n7067), .ZN(n7066) );
  OAI21_X1 U7853 ( .B1(n7068), .B2(n7070), .A(n11454), .ZN(n7067) );
  NAND2_X1 U7854 ( .A1(n6794), .A2(n7073), .ZN(n6793) );
  OR2_X1 U7855 ( .A1(n7075), .A2(n7074), .ZN(n6794) );
  NAND2_X1 U7856 ( .A1(n14358), .A2(n11453), .ZN(n7075) );
  NAND2_X1 U7857 ( .A1(n14586), .A2(n14392), .ZN(n7248) );
  AND2_X1 U7858 ( .A1(n11441), .A2(n11453), .ZN(n14359) );
  OR2_X1 U7859 ( .A1(n14372), .A2(n14373), .ZN(n7249) );
  XNOR2_X1 U7860 ( .A(n14586), .B(n14392), .ZN(n14373) );
  NAND2_X1 U7861 ( .A1(n14419), .A2(n6782), .ZN(n14400) );
  AND2_X1 U7862 ( .A1(n14413), .A2(n11451), .ZN(n14387) );
  NOR2_X1 U7863 ( .A1(n14444), .A2(n7257), .ZN(n7256) );
  INV_X1 U7864 ( .A(n11390), .ZN(n7257) );
  AOI21_X1 U7865 ( .B1(n6780), .B2(n14444), .A(n6500), .ZN(n6779) );
  INV_X1 U7866 ( .A(n11447), .ZN(n6780) );
  AOI21_X1 U7867 ( .B1(n6426), .B2(n6436), .A(n6499), .ZN(n6783) );
  AOI21_X1 U7868 ( .B1(n7266), .B2(n11350), .A(n6506), .ZN(n7265) );
  NAND2_X1 U7869 ( .A1(n11445), .A2(n12041), .ZN(n14495) );
  OR2_X1 U7870 ( .A1(n14653), .A2(n14113), .ZN(n12024) );
  OR2_X1 U7871 ( .A1(n14535), .A2(n11181), .ZN(n6789) );
  NAND2_X1 U7872 ( .A1(n6789), .A2(n6787), .ZN(n11444) );
  OAI21_X1 U7873 ( .B1(n11184), .B2(n7092), .A(n12022), .ZN(n14535) );
  INV_X1 U7874 ( .A(n12020), .ZN(n7092) );
  OR2_X1 U7875 ( .A1(n14725), .A2(n14726), .ZN(n14722) );
  NAND2_X1 U7876 ( .A1(n10530), .A2(n10529), .ZN(n14806) );
  OR2_X1 U7877 ( .A1(n10527), .A2(n9924), .ZN(n10530) );
  NOR2_X1 U7878 ( .A1(n10545), .A2(n6791), .ZN(n6790) );
  INV_X1 U7879 ( .A(n10391), .ZN(n6791) );
  OR2_X1 U7880 ( .A1(n8807), .A2(n6699), .ZN(n9271) );
  NAND2_X1 U7881 ( .A1(n7087), .A2(n7086), .ZN(n10017) );
  OR2_X1 U7882 ( .A1(n11366), .A2(n6798), .ZN(n6797) );
  NAND2_X1 U7883 ( .A1(n11907), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6798) );
  OR2_X1 U7884 ( .A1(n11391), .A2(n9219), .ZN(n9220) );
  AND2_X1 U7885 ( .A1(n9003), .A2(n9002), .ZN(n14394) );
  OR2_X1 U7886 ( .A1(n11793), .A2(n8783), .ZN(n9268) );
  AOI21_X1 U7887 ( .B1(n7074), .B2(n14343), .A(n14342), .ZN(n14575) );
  INV_X1 U7888 ( .A(n6665), .ZN(n7244) );
  OR2_X1 U7889 ( .A1(n11927), .A2(n9002), .ZN(n14637) );
  AND2_X1 U7890 ( .A1(n11171), .A2(n11170), .ZN(n14647) );
  AND2_X1 U7891 ( .A1(n11164), .A2(n14690), .ZN(n8778) );
  INV_X1 U7892 ( .A(n14135), .ZN(n14938) );
  INV_X1 U7893 ( .A(n14961), .ZN(n14949) );
  INV_X1 U7894 ( .A(n14637), .ZN(n14921) );
  INV_X1 U7895 ( .A(n14969), .ZN(n14927) );
  NAND3_X1 U7896 ( .A1(n8159), .A2(n8158), .A3(n9419), .ZN(n8163) );
  NOR2_X1 U7897 ( .A1(n8162), .A2(n7375), .ZN(n7077) );
  NAND2_X1 U7898 ( .A1(n7377), .A2(n8326), .ZN(n7375) );
  OAI21_X1 U7899 ( .B1(n11331), .B2(n7334), .A(n7333), .ZN(n11294) );
  INV_X1 U7900 ( .A(n7335), .ZN(n7334) );
  XNOR2_X1 U7901 ( .A(n8183), .B(P1_IR_REG_26__SCAN_IN), .ZN(n8347) );
  CLKBUF_X1 U7902 ( .A(n8325), .Z(n8182) );
  OAI21_X1 U7903 ( .B1(n8184), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8170) );
  NOR2_X1 U7904 ( .A1(n8763), .A2(n8172), .ZN(n8174) );
  OAI21_X1 U7905 ( .B1(n10186), .B2(n6934), .A(n6933), .ZN(n10742) );
  AND2_X1 U7906 ( .A1(n10444), .A2(n10191), .ZN(n11511) );
  NAND2_X1 U7907 ( .A1(n6514), .A2(n10443), .ZN(n10444) );
  NAND2_X1 U7908 ( .A1(n8167), .A2(n8166), .ZN(n8763) );
  OR2_X1 U7909 ( .A1(n9425), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n9534) );
  XNOR2_X1 U7910 ( .A(n8834), .B(n8833), .ZN(n10532) );
  INV_X1 U7911 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7483) );
  INV_X1 U7912 ( .A(n7481), .ZN(n7482) );
  XNOR2_X1 U7913 ( .A(n7480), .B(n7482), .ZN(n7484) );
  NOR2_X1 U7914 ( .A1(n15243), .A2(n7488), .ZN(n7490) );
  OAI21_X1 U7915 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n7454), .A(n7453), .ZN(
        n7512) );
  NAND2_X1 U7916 ( .A1(n7985), .A2(n7984), .ZN(n13155) );
  NOR2_X1 U7917 ( .A1(n9821), .A2(n7416), .ZN(n9819) );
  AOI21_X1 U7918 ( .B1(n7284), .B2(n7286), .A(n7281), .ZN(n7280) );
  INV_X1 U7919 ( .A(n12726), .ZN(n7281) );
  OR2_X1 U7920 ( .A1(n10260), .A2(n12975), .ZN(n10261) );
  AND4_X1 U7921 ( .A1(n7877), .A2(n7876), .A3(n7875), .A4(n7874), .ZN(n14775)
         );
  INV_X1 U7922 ( .A(n13221), .ZN(n13248) );
  XNOR2_X1 U7923 ( .A(n10158), .B(n9984), .ZN(n9964) );
  OAI22_X1 U7924 ( .A1(n10504), .A2(n10503), .B1(n10502), .B2(n10508), .ZN(
        n10769) );
  NAND2_X1 U7925 ( .A1(n6589), .A2(n6588), .ZN(n6587) );
  NAND2_X1 U7926 ( .A1(n11668), .A2(n7407), .ZN(n11894) );
  NAND2_X1 U7927 ( .A1(n7663), .A2(n7662), .ZN(n13309) );
  NAND2_X1 U7928 ( .A1(n7605), .A2(n7604), .ZN(n8044) );
  MUX2_X1 U7929 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7602), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n7605) );
  AND2_X1 U7930 ( .A1(n11705), .A2(n10713), .ZN(n6759) );
  XNOR2_X1 U7931 ( .A(n11723), .B(n11721), .ZN(n13437) );
  XNOR2_X1 U7932 ( .A(n9703), .B(n9704), .ZN(n9758) );
  NAND2_X1 U7933 ( .A1(n11579), .A2(n11578), .ZN(n13964) );
  NAND2_X1 U7934 ( .A1(n11104), .A2(n11069), .ZN(n11072) );
  INV_X1 U7935 ( .A(n12185), .ZN(n9834) );
  NAND2_X1 U7936 ( .A1(n11540), .A2(n11539), .ZN(n13846) );
  NAND2_X1 U7937 ( .A1(n9108), .A2(n9604), .ZN(n9609) );
  INV_X1 U7938 ( .A(n13478), .ZN(n13527) );
  NAND2_X1 U7939 ( .A1(n10684), .A2(n10683), .ZN(n12300) );
  XNOR2_X1 U7940 ( .A(n10624), .B(n10623), .ZN(n10458) );
  AND2_X1 U7941 ( .A1(n13570), .A2(n14993), .ZN(n6645) );
  XNOR2_X1 U7942 ( .A(n11646), .B(n7007), .ZN(n13947) );
  NAND2_X1 U7943 ( .A1(n11624), .A2(n11623), .ZN(n11625) );
  NAND2_X1 U7944 ( .A1(n11591), .A2(n11590), .ZN(n13954) );
  AND3_X1 U7945 ( .A1(n13830), .A2(n9326), .A3(n13829), .ZN(n13979) );
  OR2_X1 U7946 ( .A1(n8848), .A2(n8969), .ZN(n8671) );
  NAND2_X1 U7947 ( .A1(n12402), .A2(n12401), .ZN(n13940) );
  OR2_X1 U7948 ( .A1(n14074), .A2(n12399), .ZN(n12402) );
  NAND2_X1 U7949 ( .A1(n8990), .A2(n6773), .ZN(n8845) );
  INV_X1 U7950 ( .A(n12399), .ZN(n6773) );
  NAND2_X1 U7951 ( .A1(n8584), .A2(n8583), .ZN(n15084) );
  NOR2_X1 U7952 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n7384) );
  INV_X1 U7953 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8576) );
  NOR2_X1 U7954 ( .A1(n14130), .A2(n6821), .ZN(n7378) );
  INV_X1 U7955 ( .A(n9215), .ZN(n6821) );
  NOR2_X1 U7956 ( .A1(n6835), .A2(n11885), .ZN(n6834) );
  INV_X1 U7957 ( .A(n6842), .ZN(n6835) );
  NAND2_X1 U7958 ( .A1(n8967), .A2(n8966), .ZN(n9009) );
  OR2_X1 U7959 ( .A1(n8965), .A2(n11793), .ZN(n8966) );
  NAND2_X1 U7960 ( .A1(n14824), .A2(n11026), .ZN(n11031) );
  NAND2_X1 U7961 ( .A1(n10382), .A2(n10381), .ZN(n14962) );
  NAND2_X1 U7962 ( .A1(n11208), .A2(n6475), .ZN(n11215) );
  NAND2_X1 U7963 ( .A1(n14696), .A2(n11404), .ZN(n14606) );
  INV_X1 U7964 ( .A(n7106), .ZN(n7101) );
  OR2_X1 U7965 ( .A1(n11921), .A2(n9230), .ZN(n9236) );
  NAND2_X1 U7966 ( .A1(n14458), .A2(n11390), .ZN(n14445) );
  NAND2_X1 U7967 ( .A1(n14456), .A2(n11447), .ZN(n14440) );
  NAND2_X1 U7968 ( .A1(n8805), .A2(n8804), .ZN(n14541) );
  OAI21_X1 U7969 ( .B1(n14565), .B2(n14969), .A(n6945), .ZN(n14659) );
  NAND2_X1 U7970 ( .A1(n14562), .A2(n14561), .ZN(n14563) );
  AND2_X1 U7971 ( .A1(n14564), .A2(n14832), .ZN(n6946) );
  INV_X1 U7972 ( .A(n14975), .ZN(n14977) );
  INV_X1 U7973 ( .A(n7376), .ZN(n7374) );
  NAND2_X1 U7974 ( .A1(n8320), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U7975 ( .A1(n6730), .A2(n6729), .ZN(n6728) );
  NAND2_X1 U7976 ( .A1(n6736), .A2(n7506), .ZN(n6735) );
  INV_X1 U7977 ( .A(n7505), .ZN(n6736) );
  OR2_X1 U7978 ( .A1(n14853), .A2(n14852), .ZN(n6748) );
  NAND2_X1 U7979 ( .A1(n6733), .A2(n6732), .ZN(n14862) );
  INV_X1 U7980 ( .A(n7518), .ZN(n6732) );
  OAI22_X1 U7981 ( .A1(n6746), .A2(P2_ADDR_REG_18__SCAN_IN), .B1(n6747), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n6745) );
  AOI21_X1 U7982 ( .B1(n6743), .B2(n6742), .A(n6741), .ZN(n6740) );
  NAND2_X1 U7983 ( .A1(n6747), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n6742) );
  NOR3_X1 U7984 ( .A1(n6746), .A2(P2_ADDR_REG_18__SCAN_IN), .A3(n6747), .ZN(
        n6741) );
  AND2_X1 U7985 ( .A1(n11954), .A2(n12119), .ZN(n11958) );
  INV_X1 U7986 ( .A(n12217), .ZN(n6678) );
  INV_X1 U7987 ( .A(n12220), .ZN(n6671) );
  INV_X1 U7988 ( .A(n12221), .ZN(n6595) );
  INV_X1 U7989 ( .A(n11975), .ZN(n7125) );
  NAND2_X1 U7990 ( .A1(n11985), .A2(n7130), .ZN(n7129) );
  NAND2_X1 U7991 ( .A1(n7131), .A2(n11987), .ZN(n7130) );
  INV_X1 U7992 ( .A(n12249), .ZN(n6684) );
  NAND2_X1 U7993 ( .A1(n11996), .A2(n7118), .ZN(n7117) );
  INV_X1 U7994 ( .A(n11997), .ZN(n7118) );
  OAI21_X1 U7995 ( .B1(n12270), .B2(n7396), .A(n6609), .ZN(n7426) );
  AND2_X1 U7996 ( .A1(n6520), .A2(n7395), .ZN(n6609) );
  NAND2_X1 U7997 ( .A1(n12291), .A2(n6479), .ZN(n7401) );
  INV_X1 U7998 ( .A(n12295), .ZN(n6573) );
  AOI21_X1 U7999 ( .B1(n7141), .B2(n12041), .A(n7140), .ZN(n7139) );
  INV_X1 U8000 ( .A(n12040), .ZN(n7140) );
  AND2_X1 U8001 ( .A1(n12044), .A2(n7137), .ZN(n7136) );
  OR2_X1 U8002 ( .A1(n7141), .A2(n12042), .ZN(n7137) );
  AOI22_X1 U8003 ( .A1(n12300), .A2(n12408), .B1(n13547), .B2(n12403), .ZN(
        n12301) );
  NAND2_X1 U8004 ( .A1(n12055), .A2(n12057), .ZN(n7128) );
  INV_X1 U8005 ( .A(n12066), .ZN(n7134) );
  NAND2_X1 U8006 ( .A1(n6674), .A2(n6673), .ZN(n7403) );
  INV_X1 U8007 ( .A(n12317), .ZN(n6673) );
  NAND2_X1 U8008 ( .A1(n6634), .A2(n6633), .ZN(n6669) );
  INV_X1 U8009 ( .A(n12338), .ZN(n6633) );
  NAND2_X1 U8010 ( .A1(n12085), .A2(n12087), .ZN(n7120) );
  INV_X1 U8011 ( .A(n12348), .ZN(n6618) );
  INV_X1 U8012 ( .A(n12432), .ZN(n12223) );
  NAND2_X1 U8013 ( .A1(n7110), .A2(n12121), .ZN(n11933) );
  NAND2_X1 U8014 ( .A1(n7111), .A2(n11930), .ZN(n7110) );
  NAND2_X1 U8015 ( .A1(n11931), .A2(n7112), .ZN(n12121) );
  AND2_X1 U8016 ( .A1(n7018), .A2(n6471), .ZN(n7015) );
  INV_X1 U8017 ( .A(n7025), .ZN(n7024) );
  OAI21_X1 U8018 ( .B1(n7795), .B2(n7026), .A(n12932), .ZN(n7025) );
  INV_X1 U8019 ( .A(n8051), .ZN(n7026) );
  AND2_X1 U8020 ( .A1(n6766), .A2(n11692), .ZN(n6765) );
  NAND2_X1 U8021 ( .A1(n6763), .A2(n6762), .ZN(n6761) );
  INV_X1 U8022 ( .A(n13471), .ZN(n6762) );
  OR2_X1 U8023 ( .A1(n13489), .A2(n6764), .ZN(n6763) );
  CLKBUF_X3 U8024 ( .A(n12223), .Z(n12408) );
  AND2_X1 U8025 ( .A1(n6931), .A2(n6933), .ZN(n6930) );
  INV_X1 U8026 ( .A(n10741), .ZN(n6931) );
  INV_X1 U8027 ( .A(n12098), .ZN(n7116) );
  INV_X1 U8028 ( .A(n11453), .ZN(n7072) );
  AOI21_X1 U8029 ( .B1(n6920), .B2(n6922), .A(n6917), .ZN(n6916) );
  OAI21_X1 U8030 ( .B1(n6924), .B2(n11157), .A(n6926), .ZN(n6917) );
  INV_X1 U8031 ( .A(n11160), .ZN(n6926) );
  INV_X1 U8032 ( .A(n8832), .ZN(n6942) );
  OAI21_X1 U8033 ( .B1(n8968), .B2(n6771), .A(n6770), .ZN(n8258) );
  NAND2_X1 U8034 ( .A1(n6943), .A2(SI_4_), .ZN(n8256) );
  INV_X1 U8035 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7312) );
  NAND2_X1 U8036 ( .A1(n7425), .A2(n8205), .ZN(n8206) );
  INV_X1 U8037 ( .A(n8236), .ZN(n6602) );
  INV_X1 U8038 ( .A(n13125), .ZN(n12565) );
  AND2_X1 U8039 ( .A1(n12716), .A2(n7291), .ZN(n7290) );
  OR2_X1 U8040 ( .A1(n12641), .A2(n7292), .ZN(n7291) );
  INV_X1 U8041 ( .A(n12563), .ZN(n7292) );
  NAND2_X1 U8042 ( .A1(n12918), .A2(n12912), .ZN(n12952) );
  NOR2_X1 U8043 ( .A1(n12950), .A2(n12951), .ZN(n7166) );
  INV_X1 U8044 ( .A(n12952), .ZN(n7167) );
  NAND2_X1 U8045 ( .A1(n9178), .A2(n9199), .ZN(n9180) );
  AOI22_X1 U8046 ( .A1(n13021), .A2(n13020), .B1(P3_REG1_REG_16__SCAN_IN), 
        .B2(n13029), .ZN(n13046) );
  OR2_X1 U8047 ( .A1(n11669), .A2(n13089), .ZN(n12914) );
  AND2_X1 U8048 ( .A1(n11669), .A2(n13089), .ZN(n12920) );
  INV_X1 U8049 ( .A(n13109), .ZN(n13106) );
  NAND2_X1 U8050 ( .A1(n7626), .A2(n13689), .ZN(n7986) );
  INV_X1 U8051 ( .A(n7977), .ZN(n7626) );
  INV_X1 U8052 ( .A(n13225), .ZN(n7045) );
  OR2_X1 U8053 ( .A1(n6873), .A2(n6874), .ZN(n6870) );
  OR2_X1 U8054 ( .A1(n7902), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7917) );
  AND2_X1 U8055 ( .A1(n12812), .A2(n12811), .ZN(n12932) );
  INV_X1 U8056 ( .A(n11650), .ZN(n7176) );
  NAND2_X1 U8057 ( .A1(n6913), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7607) );
  INV_X1 U8058 ( .A(n7584), .ZN(n7171) );
  AND2_X1 U8059 ( .A1(n6432), .A2(n6502), .ZN(n7310) );
  INV_X1 U8060 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7600) );
  AND4_X1 U8061 ( .A1(n7598), .A2(n7597), .A3(n7596), .A4(n7656), .ZN(n7415)
         );
  INV_X1 U8062 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7596) );
  NOR2_X1 U8063 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n7598) );
  NOR2_X1 U8064 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n7597) );
  INV_X1 U8065 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7657) );
  NAND2_X1 U8066 ( .A1(n9749), .A2(n9698), .ZN(n9747) );
  OR2_X1 U8067 ( .A1(n13516), .A2(n13420), .ZN(n7239) );
  AND2_X1 U8068 ( .A1(n12380), .A2(n12381), .ZN(n6687) );
  NOR2_X1 U8069 ( .A1(n12418), .A2(n12417), .ZN(n12419) );
  NAND2_X1 U8070 ( .A1(n10946), .A2(n6957), .ZN(n6956) );
  INV_X1 U8071 ( .A(n6958), .ZN(n6957) );
  NAND2_X1 U8072 ( .A1(n10919), .A2(n6959), .ZN(n6958) );
  AND2_X1 U8073 ( .A1(n6463), .A2(n6994), .ZN(n6990) );
  INV_X1 U8074 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9488) );
  INV_X1 U8075 ( .A(n12458), .ZN(n6977) );
  NOR2_X1 U8076 ( .A1(n13414), .A2(n9750), .ZN(n7210) );
  NAND2_X1 U8077 ( .A1(n13414), .A2(n9750), .ZN(n7211) );
  NOR2_X1 U8078 ( .A1(n7209), .A2(n7210), .ZN(n7208) );
  NOR2_X1 U8079 ( .A1(n6425), .A2(n7186), .ZN(n7184) );
  INV_X1 U8080 ( .A(n11628), .ZN(n13765) );
  NAND2_X1 U8081 ( .A1(n13835), .A2(n11549), .ZN(n7206) );
  NAND2_X1 U8082 ( .A1(n10205), .A2(n10204), .ZN(n12273) );
  INV_X1 U8083 ( .A(n6951), .ZN(n9910) );
  INV_X1 U8084 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8496) );
  INV_X1 U8085 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8152) );
  OR2_X1 U8086 ( .A1(n8356), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8359) );
  INV_X1 U8087 ( .A(n11861), .ZN(n7364) );
  NOR2_X1 U8088 ( .A1(n14149), .A2(n7371), .ZN(n7370) );
  INV_X1 U8089 ( .A(n11831), .ZN(n7371) );
  INV_X1 U8090 ( .A(n11835), .ZN(n6863) );
  AOI21_X1 U8091 ( .B1(n7366), .B2(n7369), .A(n6496), .ZN(n7365) );
  INV_X1 U8092 ( .A(n11841), .ZN(n7369) );
  AND2_X1 U8093 ( .A1(n7366), .A2(n6862), .ZN(n6861) );
  OR2_X1 U8094 ( .A1(n7370), .A2(n6863), .ZN(n6862) );
  OR2_X1 U8095 ( .A1(n9229), .A2(n8390), .ZN(n8789) );
  OR2_X1 U8096 ( .A1(n11435), .A2(n8787), .ZN(n8791) );
  CLKBUF_X1 U8097 ( .A(n8635), .Z(n9420) );
  INV_X1 U8098 ( .A(n7071), .ZN(n7070) );
  OAI21_X1 U8099 ( .B1(n14359), .B2(n7072), .A(n7074), .ZN(n7071) );
  INV_X1 U8100 ( .A(n14373), .ZN(n12153) );
  INV_X1 U8101 ( .A(n11416), .ZN(n11345) );
  OR2_X1 U8102 ( .A1(n7096), .A2(n7095), .ZN(n7094) );
  INV_X1 U8103 ( .A(n6787), .ZN(n6786) );
  INV_X1 U8104 ( .A(n7088), .ZN(n7083) );
  INV_X1 U8105 ( .A(n9943), .ZN(n7085) );
  INV_X1 U8106 ( .A(n9504), .ZN(n12129) );
  AOI21_X1 U8107 ( .B1(n7247), .B2(n7246), .A(n6515), .ZN(n7245) );
  INV_X1 U8108 ( .A(n7248), .ZN(n7246) );
  NOR2_X1 U8109 ( .A1(n14501), .A2(n14489), .ZN(n6801) );
  OAI21_X1 U8110 ( .B1(n11317), .B2(n11316), .A(n11298), .ZN(n11903) );
  INV_X1 U8111 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7377) );
  AOI21_X1 U8112 ( .B1(n7335), .B2(n7337), .A(n6556), .ZN(n7333) );
  INV_X1 U8113 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8326) );
  NAND2_X1 U8114 ( .A1(n10188), .A2(SI_20_), .ZN(n6933) );
  NOR2_X1 U8115 ( .A1(n10188), .A2(SI_20_), .ZN(n6934) );
  AOI21_X1 U8116 ( .B1(n7329), .B2(n7331), .A(n7327), .ZN(n7326) );
  INV_X1 U8117 ( .A(n10184), .ZN(n7327) );
  NAND2_X1 U8118 ( .A1(n10186), .A2(n10185), .ZN(n10187) );
  INV_X1 U8119 ( .A(n10189), .ZN(n10188) );
  NAND2_X1 U8120 ( .A1(n10443), .A2(n10187), .ZN(n10190) );
  NAND2_X1 U8121 ( .A1(n6932), .A2(SI_20_), .ZN(n10443) );
  INV_X1 U8122 ( .A(n10186), .ZN(n6932) );
  NAND2_X1 U8123 ( .A1(n6563), .A2(n10082), .ZN(n10194) );
  AOI21_X1 U8124 ( .B1(n7347), .B2(n7345), .A(n9411), .ZN(n7344) );
  NAND2_X1 U8125 ( .A1(n8833), .A2(n8832), .ZN(n6941) );
  NAND2_X1 U8126 ( .A1(n8464), .A2(n8465), .ZN(n7325) );
  INV_X1 U8127 ( .A(n8466), .ZN(n8465) );
  OAI21_X1 U8128 ( .B1(n6943), .B2(SI_4_), .A(n8256), .ZN(n8243) );
  OAI21_X1 U8129 ( .B1(n8236), .B2(n9219), .A(n6661), .ZN(n8237) );
  NAND2_X1 U8130 ( .A1(n8236), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6661) );
  NAND2_X1 U8131 ( .A1(n8220), .A2(n8219), .ZN(n8233) );
  NAND2_X1 U8132 ( .A1(n8221), .A2(SI_2_), .ZN(n8235) );
  NAND2_X1 U8133 ( .A1(n8206), .A2(SI_1_), .ZN(n8232) );
  NAND2_X1 U8134 ( .A1(n6819), .A2(n7433), .ZN(n7434) );
  AOI21_X1 U8135 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n7447), .A(n7446), .ZN(
        n7448) );
  NOR2_X1 U8136 ( .A1(n7475), .A2(n7474), .ZN(n7446) );
  NAND2_X1 U8137 ( .A1(n12514), .A2(n6454), .ZN(n12591) );
  NAND2_X1 U8138 ( .A1(n12591), .A2(n12516), .ZN(n12630) );
  INV_X1 U8139 ( .A(n12526), .ZN(n7286) );
  INV_X1 U8140 ( .A(n7285), .ZN(n7284) );
  OAI21_X1 U8141 ( .B1(n12573), .B2(n7286), .A(n12725), .ZN(n7285) );
  OR2_X1 U8142 ( .A1(n7986), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7996) );
  INV_X1 U8143 ( .A(n15172), .ZN(n10093) );
  INV_X1 U8144 ( .A(n7962), .ZN(n7625) );
  INV_X1 U8145 ( .A(n7301), .ZN(n7300) );
  AOI21_X1 U8146 ( .B1(n7301), .B2(n7299), .A(n6478), .ZN(n7298) );
  NOR2_X1 U8147 ( .A1(n10674), .A2(n7294), .ZN(n7293) );
  INV_X1 U8148 ( .A(n10613), .ZN(n7294) );
  OR2_X1 U8149 ( .A1(n7767), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7780) );
  INV_X1 U8150 ( .A(n12719), .ZN(n12731) );
  OR2_X1 U8151 ( .A1(n12525), .A2(n13247), .ZN(n12526) );
  OR2_X1 U8152 ( .A1(n8122), .A2(n8121), .ZN(n9787) );
  NAND2_X1 U8153 ( .A1(n7852), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7713) );
  OR2_X1 U8154 ( .A1(n9285), .A2(n9161), .ZN(n9286) );
  NAND2_X1 U8155 ( .A1(n6585), .A2(n6584), .ZN(n9152) );
  OR2_X1 U8156 ( .A1(n13037), .A2(n9174), .ZN(n6585) );
  NAND2_X1 U8157 ( .A1(n13037), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n6584) );
  NAND2_X1 U8158 ( .A1(n9286), .A2(n9162), .ZN(n9196) );
  NAND2_X1 U8159 ( .A1(n9200), .A2(n9201), .ZN(n9199) );
  NOR2_X1 U8160 ( .A1(n15118), .A2(n15119), .ZN(n15117) );
  XNOR2_X1 U8161 ( .A(n10163), .B(n9984), .ZN(n9971) );
  NAND2_X1 U8162 ( .A1(n9971), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n10165) );
  OAI21_X1 U8163 ( .B1(n15125), .B2(n9989), .A(n9988), .ZN(n10153) );
  XNOR2_X1 U8164 ( .A(n10342), .B(n7847), .ZN(n10169) );
  NAND2_X1 U8165 ( .A1(n10169), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n10344) );
  NAND2_X1 U8166 ( .A1(n11273), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n13002) );
  INV_X1 U8167 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n13069) );
  AND2_X1 U8168 ( .A1(n13042), .A2(n6756), .ZN(n13060) );
  NAND2_X1 U8169 ( .A1(n13043), .A2(n13044), .ZN(n6756) );
  NOR2_X1 U8170 ( .A1(n13038), .A2(n6580), .ZN(n13055) );
  NOR2_X1 U8171 ( .A1(n6582), .A2(n6581), .ZN(n6580) );
  INV_X1 U8172 ( .A(n13039), .ZN(n6582) );
  NAND2_X1 U8173 ( .A1(n12903), .A2(n12904), .ZN(n7043) );
  NAND2_X1 U8174 ( .A1(n6718), .A2(n8026), .ZN(n8028) );
  NAND2_X1 U8175 ( .A1(n13108), .A2(n8025), .ZN(n6718) );
  OR2_X1 U8176 ( .A1(n8020), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8038) );
  AND2_X1 U8177 ( .A1(n12893), .A2(n12894), .ZN(n13109) );
  INV_X1 U8178 ( .A(n13135), .ZN(n13110) );
  NAND2_X1 U8179 ( .A1(n6881), .A2(n6880), .ZN(n13149) );
  AOI21_X1 U8180 ( .B1(n6885), .B2(n6879), .A(n6511), .ZN(n6883) );
  NAND2_X1 U8181 ( .A1(n7623), .A2(n7622), .ZN(n7673) );
  OR2_X1 U8182 ( .A1(n6899), .A2(n6460), .ZN(n6896) );
  NOR2_X1 U8183 ( .A1(n6460), .A2(n6898), .ZN(n6897) );
  INV_X1 U8184 ( .A(n13266), .ZN(n13260) );
  NOR2_X1 U8185 ( .A1(n7871), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7872) );
  INV_X1 U8186 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n7686) );
  AND2_X1 U8187 ( .A1(n12837), .A2(n7035), .ZN(n14758) );
  INV_X1 U8188 ( .A(n12938), .ZN(n11096) );
  OR2_X1 U8189 ( .A1(n7833), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7853) );
  OR2_X1 U8190 ( .A1(n7853), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7871) );
  INV_X1 U8191 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n7830) );
  NAND2_X1 U8192 ( .A1(n6912), .A2(n6907), .ZN(n10817) );
  NOR2_X1 U8193 ( .A1(n7797), .A2(n6908), .ZN(n6907) );
  INV_X1 U8194 ( .A(n7888), .ZN(n6908) );
  NOR2_X1 U8195 ( .A1(n7780), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7800) );
  AND2_X1 U8196 ( .A1(n7800), .A2(n7799), .ZN(n7831) );
  NAND2_X1 U8197 ( .A1(n10597), .A2(n7795), .ZN(n10596) );
  NAND2_X1 U8198 ( .A1(n10447), .A2(n12928), .ZN(n10446) );
  AND2_X1 U8199 ( .A1(n12800), .A2(n12799), .ZN(n12928) );
  AND2_X1 U8200 ( .A1(n12793), .A2(n12798), .ZN(n12931) );
  OR2_X1 U8201 ( .A1(n10576), .A2(n12931), .ZN(n10578) );
  AND2_X1 U8202 ( .A1(n8066), .A2(n8110), .ZN(n15177) );
  NOR2_X1 U8203 ( .A1(n9672), .A2(n15226), .ZN(n9800) );
  OAI21_X1 U8204 ( .B1(n15189), .B2(n9822), .A(n7710), .ZN(n15171) );
  NAND2_X1 U8205 ( .A1(n8017), .A2(n8016), .ZN(n12564) );
  NAND2_X1 U8206 ( .A1(n8116), .A2(n8120), .ZN(n9671) );
  CLKBUF_X1 U8207 ( .A(n9774), .Z(n8089) );
  NAND2_X1 U8208 ( .A1(n7582), .A2(n7583), .ZN(n7994) );
  XNOR2_X1 U8209 ( .A(n8105), .B(n8104), .ZN(n9660) );
  NAND2_X1 U8210 ( .A1(n8103), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8105) );
  INV_X1 U8211 ( .A(n7181), .ZN(n7180) );
  AOI21_X1 U8212 ( .B1(n7179), .B2(n7181), .A(n6554), .ZN(n7178) );
  NOR2_X1 U8213 ( .A1(n7641), .A2(n7182), .ZN(n7181) );
  NAND2_X1 U8214 ( .A1(n7667), .A2(n7572), .ZN(n7651) );
  AND2_X1 U8215 ( .A1(n7574), .A2(n7573), .ZN(n7650) );
  INV_X1 U8216 ( .A(n7659), .ZN(n7944) );
  AND2_X1 U8217 ( .A1(n7559), .A2(n7558), .ZN(n7882) );
  AND2_X1 U8218 ( .A1(n7555), .A2(n7554), .ZN(n7824) );
  AND2_X1 U8219 ( .A1(n7553), .A2(n7552), .ZN(n7841) );
  INV_X1 U8220 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7807) );
  OR2_X1 U8221 ( .A1(n7806), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n7809) );
  OR2_X1 U8222 ( .A1(n7809), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7838) );
  INV_X1 U8223 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7786) );
  AND2_X1 U8224 ( .A1(n7540), .A2(n7539), .ZN(n7732) );
  OR2_X1 U8225 ( .A1(n9489), .A2(n9488), .ZN(n9709) );
  AND2_X1 U8226 ( .A1(n11686), .A2(n13490), .ZN(n6766) );
  AOI21_X1 U8227 ( .B1(n10207), .B2(n9854), .A(n6449), .ZN(n7229) );
  OR2_X1 U8228 ( .A1(n11580), .A2(n13727), .ZN(n11582) );
  NAND2_X1 U8229 ( .A1(n10685), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n10934) );
  OR2_X1 U8230 ( .A1(n11233), .A2(n11232), .ZN(n11516) );
  NAND2_X1 U8231 ( .A1(n11476), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n11542) );
  INV_X1 U8232 ( .A(n11516), .ZN(n11476) );
  XNOR2_X1 U8233 ( .A(n12273), .B(n6627), .ZN(n10230) );
  AND2_X1 U8234 ( .A1(n11680), .A2(n11674), .ZN(n7233) );
  AND2_X1 U8235 ( .A1(n12498), .A2(n12441), .ZN(n9117) );
  NAND2_X1 U8236 ( .A1(n8491), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8492) );
  NAND2_X1 U8237 ( .A1(n14989), .A2(n14990), .ZN(n14988) );
  NAND2_X1 U8238 ( .A1(n15004), .A2(n15005), .ZN(n15002) );
  NAND2_X1 U8239 ( .A1(n8585), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6947) );
  NAND2_X1 U8240 ( .A1(n15017), .A2(n15018), .ZN(n15016) );
  AND2_X1 U8241 ( .A1(n8537), .A2(n8538), .ZN(n8535) );
  AOI21_X1 U8242 ( .B1(n9483), .B2(P2_REG2_REG_8__SCAN_IN), .A(n15037), .ZN(
        n8519) );
  AOI21_X1 U8243 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n9841), .A(n8890), .ZN(
        n8893) );
  AOI21_X1 U8244 ( .B1(n10203), .B2(P2_REG1_REG_11__SCAN_IN), .A(n9064), .ZN(
        n9065) );
  NAND2_X1 U8245 ( .A1(n9068), .A2(n6590), .ZN(n9069) );
  OR2_X1 U8246 ( .A1(n10203), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6590) );
  NAND2_X1 U8247 ( .A1(n9069), .A2(n9070), .ZN(n9897) );
  AOI21_X1 U8248 ( .B1(n15051), .B2(P2_REG2_REG_13__SCAN_IN), .A(n15053), .ZN(
        n10461) );
  INV_X1 U8249 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11706) );
  AND2_X1 U8250 ( .A1(n6641), .A2(n6640), .ZN(n9902) );
  NAND2_X1 U8251 ( .A1(n15051), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6640) );
  NAND2_X1 U8252 ( .A1(n10630), .A2(n10631), .ZN(n10634) );
  NOR2_X1 U8253 ( .A1(n11255), .A2(n6647), .ZN(n11257) );
  AND2_X1 U8254 ( .A1(n11256), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6647) );
  AND2_X1 U8255 ( .A1(n11251), .A2(n11250), .ZN(n11253) );
  INV_X1 U8256 ( .A(n6971), .ZN(n6970) );
  INV_X1 U8257 ( .A(n6969), .ZN(n6968) );
  OAI21_X1 U8258 ( .B1(n6972), .B2(n6970), .A(n13769), .ZN(n6969) );
  NOR2_X1 U8259 ( .A1(n13960), .A2(n6953), .ZN(n6952) );
  INV_X1 U8260 ( .A(n6954), .ZN(n6953) );
  NAND2_X1 U8261 ( .A1(n11627), .A2(n13815), .ZN(n13809) );
  NAND2_X1 U8262 ( .A1(n11627), .A2(n6954), .ZN(n13794) );
  AOI21_X1 U8263 ( .B1(n6983), .B2(n6981), .A(n6490), .ZN(n6980) );
  INV_X1 U8264 ( .A(n6983), .ZN(n6982) );
  INV_X1 U8265 ( .A(n11639), .ZN(n6981) );
  NAND2_X1 U8266 ( .A1(n7200), .A2(n7198), .ZN(n13805) );
  AOI21_X1 U8267 ( .B1(n7201), .B2(n7205), .A(n7199), .ZN(n7198) );
  AOI21_X1 U8268 ( .B1(n7204), .B2(n7203), .A(n7202), .ZN(n7201) );
  NAND2_X1 U8269 ( .A1(n7206), .A2(n7204), .ZN(n13818) );
  NAND2_X1 U8270 ( .A1(n6998), .A2(n6996), .ZN(n13878) );
  AOI21_X1 U8271 ( .B1(n6451), .B2(n11633), .A(n6997), .ZN(n6996) );
  INV_X1 U8272 ( .A(n11636), .ZN(n6997) );
  NAND2_X1 U8273 ( .A1(n13890), .A2(n13896), .ZN(n13889) );
  AOI21_X1 U8274 ( .B1(n11142), .B2(n7223), .A(n6476), .ZN(n11231) );
  NOR2_X1 U8275 ( .A1(n11228), .A2(n7224), .ZN(n7223) );
  INV_X1 U8276 ( .A(n11141), .ZN(n7224) );
  NAND2_X1 U8277 ( .A1(n7002), .A2(n7001), .ZN(n11222) );
  AOI21_X1 U8278 ( .B1(n7003), .B2(n10920), .A(n6465), .ZN(n7001) );
  NOR2_X1 U8279 ( .A1(n10662), .A2(n6956), .ZN(n11147) );
  NOR2_X1 U8280 ( .A1(n10662), .A2(n6958), .ZN(n10943) );
  NOR2_X1 U8281 ( .A1(n10662), .A2(n6593), .ZN(n10694) );
  NAND2_X1 U8282 ( .A1(n10559), .A2(n7220), .ZN(n10652) );
  NOR2_X1 U8283 ( .A1(n10569), .A2(n7221), .ZN(n7220) );
  INV_X1 U8284 ( .A(n10558), .ZN(n7221) );
  NAND2_X1 U8285 ( .A1(n10213), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n10220) );
  INV_X1 U8286 ( .A(n10214), .ZN(n10213) );
  XNOR2_X1 U8287 ( .A(n15089), .B(n8952), .ZN(n12451) );
  MUX2_X1 U8288 ( .A(n8600), .B(n14090), .S(n8931), .Z(n12185) );
  NAND2_X1 U8289 ( .A1(n10931), .A2(n10930), .ZN(n10932) );
  NAND2_X1 U8290 ( .A1(n10650), .A2(n10649), .ZN(n12294) );
  NAND2_X1 U8291 ( .A1(n10212), .A2(n10211), .ZN(n12281) );
  NAND2_X1 U8292 ( .A1(n10830), .A2(n12393), .ZN(n10212) );
  NAND2_X1 U8293 ( .A1(n9482), .A2(n6979), .ZN(n9760) );
  NOR2_X1 U8294 ( .A1(n9124), .A2(n8581), .ZN(n8798) );
  NAND2_X1 U8295 ( .A1(n6448), .A2(n6630), .ZN(n11473) );
  NAND2_X1 U8296 ( .A1(n8574), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n6630) );
  INV_X1 U8297 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8140) );
  NOR2_X1 U8298 ( .A1(n9042), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n9407) );
  AND2_X1 U8299 ( .A1(n8264), .A2(n8263), .ZN(n8935) );
  INV_X1 U8300 ( .A(n14346), .ZN(n14103) );
  AND2_X1 U8301 ( .A1(n14222), .A2(n7363), .ZN(n7362) );
  OR2_X1 U8302 ( .A1(n14158), .A2(n7364), .ZN(n7363) );
  OR2_X1 U8303 ( .A1(n10841), .A2(n10840), .ZN(n10857) );
  NOR2_X1 U8304 ( .A1(n14111), .A2(n6856), .ZN(n6855) );
  INV_X1 U8305 ( .A(n7354), .ZN(n6856) );
  NAND2_X1 U8306 ( .A1(n11784), .A2(n7355), .ZN(n7354) );
  INV_X1 U8307 ( .A(n11786), .ZN(n7355) );
  INV_X1 U8308 ( .A(n11406), .ZN(n11417) );
  NAND2_X1 U8309 ( .A1(n11417), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11416) );
  NAND2_X1 U8310 ( .A1(n14194), .A2(n7370), .ZN(n14146) );
  NAND2_X1 U8311 ( .A1(n10538), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10841) );
  AND2_X1 U8312 ( .A1(n11172), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11186) );
  NAND2_X1 U8313 ( .A1(n6826), .A2(n6540), .ZN(n11795) );
  INV_X1 U8314 ( .A(n7353), .ZN(n6826) );
  AOI22_X1 U8315 ( .A1(n11875), .A2(n9573), .B1(n8711), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n8712) );
  OR2_X1 U8316 ( .A1(n11371), .A2(n11370), .ZN(n11380) );
  NOR2_X1 U8317 ( .A1(n11380), .A2(n14198), .ZN(n11395) );
  INV_X1 U8318 ( .A(n11394), .ZN(n11407) );
  NAND2_X1 U8319 ( .A1(n14146), .A2(n11835), .ZN(n14203) );
  NAND2_X1 U8320 ( .A1(n14203), .A2(n14204), .ZN(n14202) );
  AND2_X1 U8321 ( .A1(n10536), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10538) );
  NAND2_X1 U8322 ( .A1(n11874), .A2(n9387), .ZN(n8994) );
  AND2_X1 U8323 ( .A1(n11186), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11360) );
  NAND2_X1 U8324 ( .A1(n11360), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11371) );
  OR2_X1 U8325 ( .A1(n10857), .A2(n14112), .ZN(n10979) );
  AOI22_X1 U8326 ( .A1(n7106), .A2(n6526), .B1(n7102), .B2(n7107), .ZN(n7100)
         );
  AND2_X1 U8327 ( .A1(n10983), .A2(n10982), .ZN(n14113) );
  INV_X2 U8328 ( .A(n9229), .ZN(n11459) );
  NAND2_X1 U8329 ( .A1(n11301), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8701) );
  INV_X1 U8330 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n8721) );
  NOR2_X1 U8331 ( .A1(n14331), .A2(n6804), .ZN(n6803) );
  INV_X1 U8332 ( .A(n6805), .ZN(n6804) );
  NOR2_X1 U8333 ( .A1(n14572), .A2(n14243), .ZN(n6944) );
  NAND2_X1 U8334 ( .A1(n14360), .A2(n14359), .ZN(n14358) );
  INV_X1 U8335 ( .A(n11457), .ZN(n14374) );
  NAND2_X1 U8336 ( .A1(n14385), .A2(n6781), .ZN(n14370) );
  NAND2_X1 U8337 ( .A1(n6782), .A2(n14244), .ZN(n6781) );
  NAND2_X1 U8338 ( .A1(n11414), .A2(n11413), .ZN(n14420) );
  AOI21_X1 U8339 ( .B1(n6776), .B2(n14439), .A(n6494), .ZN(n6774) );
  NAND2_X1 U8340 ( .A1(n14415), .A2(n14414), .ZN(n14413) );
  AOI21_X1 U8341 ( .B1(n14430), .B2(n7254), .A(n6483), .ZN(n7253) );
  INV_X1 U8342 ( .A(n11401), .ZN(n7254) );
  NAND2_X1 U8343 ( .A1(n6802), .A2(n14507), .ZN(n14501) );
  INV_X1 U8344 ( .A(n6802), .ZN(n14520) );
  NAND2_X1 U8345 ( .A1(n14513), .A2(n12039), .ZN(n14492) );
  NAND2_X1 U8346 ( .A1(n10974), .A2(n10973), .ZN(n11184) );
  INV_X1 U8347 ( .A(n12145), .ZN(n14726) );
  NAND2_X1 U8348 ( .A1(n10707), .A2(n10531), .ZN(n10851) );
  AOI21_X1 U8349 ( .B1(n7260), .B2(n12139), .A(n6492), .ZN(n7258) );
  INV_X1 U8350 ( .A(n7260), .ZN(n7259) );
  NOR2_X1 U8351 ( .A1(n10384), .A2(n10383), .ZN(n10536) );
  NAND2_X1 U8352 ( .A1(n6800), .A2(n6799), .ZN(n10705) );
  OR2_X1 U8353 ( .A1(n10117), .A2(n10116), .ZN(n10384) );
  NAND2_X1 U8354 ( .A1(n10392), .A2(n10391), .ZN(n10393) );
  NAND2_X1 U8355 ( .A1(n7087), .A2(n7090), .ZN(n10015) );
  AND2_X1 U8356 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9253) );
  NAND2_X1 U8357 ( .A1(n11957), .A2(n11954), .ZN(n9504) );
  NAND2_X1 U8358 ( .A1(n14267), .A2(n9573), .ZN(n9389) );
  AND2_X1 U8359 ( .A1(n11770), .A2(n11769), .ZN(n14567) );
  INV_X1 U8360 ( .A(n14348), .ZN(n11768) );
  NAND2_X1 U8361 ( .A1(n11177), .A2(n11176), .ZN(n14545) );
  NAND2_X1 U8362 ( .A1(n9271), .A2(n8808), .ZN(n14961) );
  AND2_X1 U8363 ( .A1(n14497), .A2(n14966), .ZN(n14969) );
  XNOR2_X1 U8364 ( .A(n11912), .B(n11911), .ZN(n14067) );
  NAND2_X1 U8365 ( .A1(n12115), .A2(n11909), .ZN(n11912) );
  INV_X1 U8366 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8691) );
  XNOR2_X1 U8367 ( .A(n8329), .B(n8326), .ZN(n14885) );
  OAI21_X1 U8368 ( .B1(n8325), .B2(P1_IR_REG_26__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8329) );
  NAND2_X1 U8369 ( .A1(n7332), .A2(n7335), .ZN(n11327) );
  NAND2_X1 U8370 ( .A1(n11331), .A2(n7339), .ZN(n7332) );
  AND2_X1 U8371 ( .A1(n11426), .A2(n11427), .ZN(n14082) );
  NAND2_X1 U8372 ( .A1(n7341), .A2(n7339), .ZN(n11427) );
  AND2_X1 U8373 ( .A1(n11288), .A2(n11162), .ZN(n11564) );
  NAND2_X1 U8374 ( .A1(n6919), .A2(n6918), .ZN(n11161) );
  NAND2_X1 U8375 ( .A1(n6914), .A2(n6923), .ZN(n6919) );
  INV_X1 U8376 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8185) );
  AND2_X1 U8377 ( .A1(n6472), .A2(n8323), .ZN(n7135) );
  NAND2_X1 U8378 ( .A1(n8763), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8703) );
  OR2_X1 U8379 ( .A1(n9534), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n10084) );
  NAND2_X1 U8380 ( .A1(n7349), .A2(n9031), .ZN(n9037) );
  NAND2_X1 U8381 ( .A1(n8463), .A2(n8462), .ZN(n6767) );
  INV_X1 U8382 ( .A(n7325), .ZN(n7324) );
  OAI21_X1 U8383 ( .B1(n8236), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n6691), .ZN(
        n8208) );
  NAND2_X1 U8384 ( .A1(n8236), .A2(n8598), .ZN(n6691) );
  NAND2_X1 U8385 ( .A1(n7428), .A2(n6816), .ZN(n7479) );
  NAND2_X1 U8386 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n6817), .ZN(n6816) );
  INV_X1 U8387 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6817) );
  XNOR2_X1 U8388 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n7478) );
  XNOR2_X1 U8389 ( .A(n7429), .B(n6812), .ZN(n7477) );
  INV_X1 U8390 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n6812) );
  XNOR2_X1 U8391 ( .A(n7476), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n7487) );
  INV_X1 U8392 ( .A(n7506), .ZN(n6737) );
  OAI22_X1 U8393 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n7452), .B1(n7451), .B2(
        n7472), .ZN(n7471) );
  AND2_X1 U8394 ( .A1(n6810), .A2(n6811), .ZN(n7522) );
  NAND2_X1 U8395 ( .A1(n7520), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n6810) );
  NAND2_X1 U8396 ( .A1(n14866), .A2(n14867), .ZN(n7520) );
  NOR2_X1 U8397 ( .A1(n14701), .A2(n14753), .ZN(n6746) );
  NAND2_X1 U8398 ( .A1(n8101), .A2(n8100), .ZN(n9661) );
  CLKBUF_X1 U8399 ( .A(n12574), .Z(n6690) );
  NAND2_X1 U8400 ( .A1(n12514), .A2(n12513), .ZN(n12593) );
  NAND2_X1 U8401 ( .A1(n7276), .A2(n7273), .ZN(n10059) );
  INV_X1 U8402 ( .A(n7275), .ZN(n7273) );
  AND2_X1 U8403 ( .A1(n12770), .A2(n12775), .ZN(n15189) );
  NAND2_X1 U8404 ( .A1(n12674), .A2(n12546), .ZN(n12622) );
  NAND2_X1 U8405 ( .A1(n8007), .A2(n8006), .ZN(n13128) );
  AND4_X1 U8406 ( .A1(n7922), .A2(n7921), .A3(n7920), .A4(n7919), .ZN(n13235)
         );
  OR2_X1 U8407 ( .A1(n10057), .A2(n7272), .ZN(n7271) );
  NAND2_X1 U8408 ( .A1(n7270), .A2(n7279), .ZN(n7269) );
  INV_X1 U8409 ( .A(n7279), .ZN(n7272) );
  XNOR2_X1 U8410 ( .A(n10260), .B(n6635), .ZN(n10091) );
  NAND2_X1 U8411 ( .A1(n12672), .A2(n12543), .ZN(n12674) );
  INV_X1 U8412 ( .A(n12739), .ZN(n12673) );
  INV_X1 U8413 ( .A(n7304), .ZN(n7303) );
  OAI21_X1 U8414 ( .B1(n7305), .B2(n6454), .A(n12521), .ZN(n7304) );
  NAND2_X1 U8415 ( .A1(n7306), .A2(n12516), .ZN(n7305) );
  XNOR2_X1 U8416 ( .A(n12550), .B(n12549), .ZN(n12691) );
  OR2_X1 U8417 ( .A1(n9787), .A2(n12960), .ZN(n12719) );
  INV_X1 U8418 ( .A(n12734), .ZN(n12717) );
  NAND2_X1 U8419 ( .A1(n7295), .A2(n10613), .ZN(n10673) );
  NAND2_X1 U8420 ( .A1(n7289), .A2(n12563), .ZN(n12715) );
  NAND2_X1 U8421 ( .A1(n12640), .A2(n12641), .ZN(n7289) );
  NAND2_X1 U8422 ( .A1(n7283), .A2(n12526), .ZN(n12727) );
  NAND2_X1 U8423 ( .A1(n6690), .A2(n12573), .ZN(n7283) );
  INV_X1 U8424 ( .A(n12720), .ZN(n12737) );
  AND4_X1 U8425 ( .A1(n10039), .A2(n9879), .A3(n9878), .A4(n9877), .ZN(n13081)
         );
  AND4_X1 U8426 ( .A1(n10039), .A2(n9874), .A3(n9873), .A4(n9872), .ZN(n12755)
         );
  INV_X1 U8427 ( .A(n13164), .ZN(n13136) );
  XNOR2_X1 U8428 ( .A(n9152), .B(n6583), .ZN(n9283) );
  AOI22_X1 U8429 ( .A1(n9469), .A2(n9470), .B1(n9478), .B2(n9156), .ZN(n9367)
         );
  AND2_X1 U8430 ( .A1(n7746), .A2(n7745), .ZN(n9190) );
  INV_X1 U8431 ( .A(n9962), .ZN(n15115) );
  NAND2_X1 U8432 ( .A1(n10159), .A2(n10160), .ZN(n15135) );
  XNOR2_X1 U8433 ( .A(n10336), .B(n7847), .ZN(n10162) );
  AOI22_X1 U8434 ( .A1(n10769), .A2(n10768), .B1(n10767), .B2(n10766), .ZN(
        n12979) );
  NAND2_X1 U8435 ( .A1(n11116), .A2(n11117), .ZN(n11266) );
  AOI21_X1 U8436 ( .B1(n11121), .B2(n11120), .A(n11119), .ZN(n11125) );
  NOR2_X1 U8437 ( .A1(n13008), .A2(n6613), .ZN(n13012) );
  AND2_X1 U8438 ( .A1(n13009), .A2(n13010), .ZN(n6613) );
  XNOR2_X1 U8439 ( .A(n13043), .B(n6581), .ZN(n13019) );
  NAND2_X1 U8440 ( .A1(n13019), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n13042) );
  XNOR2_X1 U8441 ( .A(n13055), .B(n13058), .ZN(n13040) );
  INV_X1 U8442 ( .A(n13277), .ZN(n13095) );
  AND2_X1 U8443 ( .A1(n7054), .A2(n12766), .ZN(n13122) );
  NAND2_X1 U8444 ( .A1(n6894), .A2(n6893), .ZN(n13123) );
  INV_X1 U8445 ( .A(n7054), .ZN(n13138) );
  NAND2_X1 U8446 ( .A1(n6882), .A2(n6885), .ZN(n13161) );
  NAND2_X1 U8447 ( .A1(n13183), .A2(n6886), .ZN(n6882) );
  OAI21_X1 U8448 ( .B1(n13189), .B2(n7018), .A(n7017), .ZN(n13166) );
  AOI21_X1 U8449 ( .B1(n13183), .B2(n12944), .A(n6428), .ZN(n13172) );
  NAND2_X1 U8450 ( .A1(n13187), .A2(n12873), .ZN(n13176) );
  NAND2_X1 U8451 ( .A1(n6900), .A2(n6901), .ZN(n13208) );
  NAND2_X1 U8452 ( .A1(n13224), .A2(n12857), .ZN(n13213) );
  AND2_X1 U8453 ( .A1(n13224), .A2(n7047), .ZN(n13212) );
  OAI21_X1 U8454 ( .B1(n14757), .B2(n7033), .A(n7030), .ZN(n13238) );
  INV_X1 U8455 ( .A(n6872), .ZN(n13245) );
  AOI21_X1 U8456 ( .B1(n6875), .B2(n6874), .A(n6873), .ZN(n6872) );
  NAND2_X1 U8457 ( .A1(n7029), .A2(n7034), .ZN(n13250) );
  NAND2_X1 U8458 ( .A1(n14757), .A2(n6453), .ZN(n7029) );
  NAND2_X1 U8459 ( .A1(n14757), .A2(n12837), .ZN(n7036) );
  NAND2_X1 U8460 ( .A1(n10880), .A2(n7052), .ZN(n14771) );
  NOR2_X1 U8461 ( .A1(n9802), .A2(n15182), .ZN(n14770) );
  INV_X1 U8462 ( .A(n15200), .ZN(n15182) );
  NAND2_X1 U8463 ( .A1(n13072), .A2(n9775), .ZN(n15200) );
  INV_X2 U8464 ( .A(n15204), .ZN(n15206) );
  NAND2_X1 U8465 ( .A1(n9802), .A2(n15169), .ZN(n15204) );
  NAND2_X1 U8466 ( .A1(n14770), .A2(n13311), .ZN(n15165) );
  NAND2_X1 U8467 ( .A1(n15240), .A2(n13311), .ZN(n13334) );
  INV_X1 U8468 ( .A(n12756), .ZN(n13337) );
  NAND2_X1 U8469 ( .A1(n12752), .A2(n12751), .ZN(n13339) );
  INV_X1 U8470 ( .A(n6708), .ZN(n6707) );
  INV_X1 U8471 ( .A(n11894), .ZN(n6710) );
  OAI21_X1 U8472 ( .B1(n11901), .B2(n14790), .A(n6709), .ZN(n6708) );
  OR2_X1 U8473 ( .A1(n13103), .A2(n8067), .ZN(n8127) );
  INV_X1 U8474 ( .A(n12899), .ZN(n13101) );
  INV_X1 U8475 ( .A(n12564), .ZN(n13348) );
  OR2_X1 U8476 ( .A1(n7749), .A2(n8273), .ZN(n7708) );
  OR2_X1 U8477 ( .A1(n15234), .A2(n15226), .ZN(n13384) );
  AND2_X1 U8478 ( .A1(n8083), .A2(n8082), .ZN(n13386) );
  AND2_X1 U8479 ( .A1(n9660), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13387) );
  XNOR2_X1 U8480 ( .A(n7152), .B(n12745), .ZN(n13394) );
  OAI21_X1 U8481 ( .B1(n12743), .B2(n12742), .A(n12744), .ZN(n7152) );
  NAND2_X1 U8482 ( .A1(n7616), .A2(n7615), .ZN(n7617) );
  NAND2_X1 U8483 ( .A1(n7610), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7615) );
  NAND2_X1 U8484 ( .A1(n7177), .A2(n11650), .ZN(n11657) );
  OR2_X1 U8485 ( .A1(n11649), .A2(n11648), .ZN(n7177) );
  INV_X1 U8486 ( .A(n8086), .ZN(n10809) );
  NAND2_X1 U8487 ( .A1(n7971), .A2(n7578), .ZN(n7642) );
  AND2_X1 U8488 ( .A1(n6772), .A2(P3_U3151), .ZN(n13393) );
  NAND2_X1 U8489 ( .A1(n8035), .A2(n8068), .ZN(n10042) );
  INV_X1 U8490 ( .A(n8117), .ZN(n9775) );
  INV_X1 U8491 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7660) );
  OAI21_X1 U8492 ( .B1(n7668), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7661) );
  INV_X1 U8493 ( .A(SI_19_), .ZN(n10198) );
  OAI21_X1 U8494 ( .B1(n7928), .B2(n7159), .A(n7156), .ZN(n7665) );
  NAND2_X1 U8495 ( .A1(n7941), .A2(n7940), .ZN(n7943) );
  NAND2_X1 U8496 ( .A1(n7928), .A2(n7568), .ZN(n7941) );
  INV_X1 U8497 ( .A(SI_16_), .ZN(n13618) );
  INV_X1 U8498 ( .A(SI_15_), .ZN(n9538) );
  OAI21_X1 U8499 ( .B1(n7680), .B2(n7164), .A(n7162), .ZN(n7910) );
  INV_X1 U8500 ( .A(SI_14_), .ZN(n9413) );
  NAND2_X1 U8501 ( .A1(n7896), .A2(n7895), .ZN(n7898) );
  NAND2_X1 U8502 ( .A1(n7680), .A2(n7562), .ZN(n7896) );
  NAND2_X1 U8503 ( .A1(n7561), .A2(n7562), .ZN(n7678) );
  INV_X1 U8504 ( .A(SI_13_), .ZN(n9033) );
  INV_X1 U8505 ( .A(SI_11_), .ZN(n8830) );
  NAND2_X1 U8506 ( .A1(n7792), .A2(n7548), .ZN(n7812) );
  NAND2_X1 U8507 ( .A1(n7146), .A2(n7147), .ZN(n7790) );
  NAND2_X1 U8508 ( .A1(n7148), .A2(n7545), .ZN(n7776) );
  NAND2_X1 U8509 ( .A1(n7762), .A2(n7761), .ZN(n7148) );
  INV_X1 U8510 ( .A(n7534), .ZN(n7699) );
  AND2_X1 U8511 ( .A1(n6441), .A2(n13427), .ZN(n7235) );
  NAND2_X1 U8512 ( .A1(n9856), .A2(n9855), .ZN(n11744) );
  NAND2_X1 U8513 ( .A1(n11490), .A2(n11489), .ZN(n13608) );
  XNOR2_X1 U8514 ( .A(n10406), .B(n10407), .ZN(n10232) );
  NAND2_X1 U8515 ( .A1(n6564), .A2(n11066), .ZN(n11106) );
  INV_X1 U8516 ( .A(n11107), .ZN(n7231) );
  AOI21_X1 U8517 ( .B1(n7243), .B2(n7241), .A(n6421), .ZN(n7240) );
  INV_X1 U8518 ( .A(n9702), .ZN(n7241) );
  OR2_X1 U8519 ( .A1(n13478), .A2(n9326), .ZN(n13512) );
  AND2_X1 U8520 ( .A1(n6424), .A2(n11686), .ZN(n13491) );
  NAND2_X1 U8521 ( .A1(n6683), .A2(n6682), .ZN(n11704) );
  INV_X1 U8522 ( .A(n10415), .ZN(n6682) );
  NAND2_X1 U8523 ( .A1(n13540), .A2(n6649), .ZN(n6648) );
  NAND2_X1 U8524 ( .A1(n11744), .A2(n10207), .ZN(n11755) );
  XNOR2_X1 U8525 ( .A(n10230), .B(n10208), .ZN(n11745) );
  NAND2_X1 U8526 ( .A1(n7228), .A2(n7227), .ZN(n9726) );
  NOR2_X1 U8527 ( .A1(n9728), .A2(n9105), .ZN(n7227) );
  NAND2_X1 U8528 ( .A1(n11675), .A2(n11674), .ZN(n13507) );
  NAND2_X1 U8529 ( .A1(n9119), .A2(n12494), .ZN(n13503) );
  NAND2_X1 U8530 ( .A1(n7234), .A2(n7236), .ZN(n13528) );
  AOI21_X1 U8531 ( .B1(n13480), .B2(n11735), .A(n11734), .ZN(n13421) );
  CLKBUF_X1 U8532 ( .A(n11067), .Z(n6564) );
  NAND2_X1 U8533 ( .A1(n11599), .A2(n11598), .ZN(n13535) );
  OR2_X1 U8534 ( .A1(n13763), .A2(n11606), .ZN(n11599) );
  NAND2_X1 U8535 ( .A1(n12390), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8609) );
  AND2_X1 U8536 ( .A1(n8607), .A2(n8608), .ZN(n6961) );
  CLKBUF_X1 U8537 ( .A(n12180), .Z(n13563) );
  OR2_X2 U8538 ( .A1(n9093), .A2(n8156), .ZN(n13562) );
  NAND2_X1 U8539 ( .A1(n15026), .A2(n15025), .ZN(n15024) );
  AOI21_X1 U8540 ( .B1(n9483), .B2(P2_REG1_REG_8__SCAN_IN), .A(n15029), .ZN(
        n8487) );
  AOI21_X1 U8541 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n9841), .A(n8884), .ZN(
        n8886) );
  INV_X1 U8542 ( .A(n6641), .ZN(n15045) );
  AND2_X1 U8543 ( .A1(n8521), .A2(n8520), .ZN(n15039) );
  NOR2_X1 U8544 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n11254), .ZN(n13567) );
  INV_X1 U8545 ( .A(n11647), .ZN(n7006) );
  NAND2_X1 U8546 ( .A1(n13949), .A2(n13808), .ZN(n13606) );
  NAND2_X1 U8547 ( .A1(n6967), .A2(n6971), .ZN(n13768) );
  NAND2_X1 U8548 ( .A1(n13792), .A2(n6972), .ZN(n6967) );
  OAI21_X1 U8549 ( .B1(n13792), .B2(n6970), .A(n6968), .ZN(n13952) );
  NAND2_X1 U8550 ( .A1(n7191), .A2(n6458), .ZN(n13759) );
  NAND2_X1 U8551 ( .A1(n13772), .A2(n7192), .ZN(n7191) );
  AND2_X1 U8552 ( .A1(n6974), .A2(n6975), .ZN(n13782) );
  NAND2_X1 U8553 ( .A1(n13792), .A2(n11643), .ZN(n6974) );
  NAND2_X1 U8554 ( .A1(n13838), .A2(n11639), .ZN(n13828) );
  NAND2_X1 U8555 ( .A1(n11553), .A2(n11552), .ZN(n13977) );
  NAND2_X1 U8556 ( .A1(n7219), .A2(n11524), .ZN(n13856) );
  NAND2_X1 U8557 ( .A1(n7000), .A2(n11635), .ZN(n13895) );
  OR2_X1 U8558 ( .A1(n11634), .A2(n11633), .ZN(n7000) );
  NAND2_X1 U8559 ( .A1(n11227), .A2(n11226), .ZN(n14006) );
  NAND2_X1 U8560 ( .A1(n11142), .A2(n11141), .ZN(n11229) );
  NAND2_X1 U8561 ( .A1(n7004), .A2(n7003), .ZN(n11145) );
  NAND2_X1 U8562 ( .A1(n7004), .A2(n10922), .ZN(n10926) );
  NAND2_X1 U8563 ( .A1(n6995), .A2(n6994), .ZN(n10698) );
  NAND2_X1 U8564 ( .A1(n6993), .A2(n6991), .ZN(n6995) );
  NAND2_X1 U8565 ( .A1(n6993), .A2(n10568), .ZN(n10661) );
  OAI21_X1 U8566 ( .B1(n9765), .B2(n7197), .A(n6430), .ZN(n9914) );
  NAND2_X1 U8567 ( .A1(n9766), .A2(n12460), .ZN(n9913) );
  NAND2_X1 U8568 ( .A1(n9765), .A2(n9764), .ZN(n9766) );
  NAND2_X1 U8569 ( .A1(n10311), .A2(n9441), .ZN(n9485) );
  INV_X1 U8570 ( .A(n13923), .ZN(n13866) );
  NAND2_X1 U8571 ( .A1(n15087), .A2(n9100), .ZN(n13825) );
  INV_X1 U8572 ( .A(n13866), .ZN(n15064) );
  NOR2_X1 U8573 ( .A1(n15075), .A2(n13603), .ZN(n13923) );
  OR2_X1 U8574 ( .A1(n10098), .A2(n12399), .ZN(n6565) );
  INV_X1 U8575 ( .A(n14015), .ZN(n13992) );
  INV_X1 U8576 ( .A(n13579), .ZN(n14024) );
  INV_X1 U8577 ( .A(n13940), .ZN(n14028) );
  AND2_X1 U8578 ( .A1(n13945), .A2(n6659), .ZN(n6658) );
  NAND2_X1 U8579 ( .A1(n6660), .A2(n14012), .ZN(n6659) );
  INV_X1 U8580 ( .A(n13608), .ZN(n14032) );
  NOR2_X1 U8581 ( .A1(n13948), .A2(n7216), .ZN(n7215) );
  NAND2_X1 U8582 ( .A1(n7217), .A2(n6485), .ZN(n7216) );
  NAND2_X1 U8583 ( .A1(n13949), .A2(n14012), .ZN(n7217) );
  NAND2_X1 U8584 ( .A1(n11527), .A2(n11526), .ZN(n14050) );
  INV_X1 U8585 ( .A(n13899), .ZN(n14059) );
  OR2_X1 U8587 ( .A1(n10527), .A2(n12399), .ZN(n9843) );
  AND2_X2 U8588 ( .A1(n8798), .A2(n15084), .ZN(n15106) );
  AND2_X1 U8589 ( .A1(n9093), .A2(n8578), .ZN(n15087) );
  NAND2_X1 U8590 ( .A1(n6963), .A2(n6962), .ZN(n8592) );
  NAND2_X1 U8591 ( .A1(n8588), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6962) );
  CLKBUF_X1 U8592 ( .A(n8500), .Z(n8501) );
  NAND2_X1 U8593 ( .A1(n8493), .A2(n8149), .ZN(n14084) );
  NAND2_X1 U8594 ( .A1(n9593), .A2(n7213), .ZN(n8147) );
  XNOR2_X1 U8595 ( .A(n8150), .B(n13732), .ZN(n14089) );
  XNOR2_X1 U8596 ( .A(n8142), .B(P2_IR_REG_24__SCAN_IN), .ZN(n11165) );
  NAND2_X1 U8597 ( .A1(n7350), .A2(n10798), .ZN(n10799) );
  INV_X1 U8598 ( .A(n7351), .ZN(n7350) );
  INV_X1 U8599 ( .A(n12441), .ZN(n12179) );
  INV_X1 U8600 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10083) );
  INV_X1 U8601 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9415) );
  INV_X1 U8602 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9080) );
  INV_X1 U8603 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n8840) );
  INV_X1 U8604 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n8633) );
  INV_X1 U8605 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n8469) );
  INV_X1 U8606 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n8382) );
  INV_X1 U8607 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n8318) );
  INV_X1 U8608 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n8285) );
  INV_X1 U8609 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n8246) );
  AND2_X1 U8610 ( .A1(n8229), .A2(n8259), .ZN(n15009) );
  INV_X1 U8611 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8850) );
  NAND2_X1 U8612 ( .A1(n8251), .A2(n8250), .ZN(n8849) );
  NAND2_X1 U8613 ( .A1(n8217), .A2(n8248), .ZN(n14992) );
  INV_X1 U8614 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8669) );
  NAND2_X1 U8615 ( .A1(n8215), .A2(n8214), .ZN(n8672) );
  NAND2_X1 U8616 ( .A1(n6846), .A2(n6850), .ZN(n14094) );
  OR2_X1 U8617 ( .A1(n9615), .A2(n6851), .ZN(n6846) );
  NAND2_X1 U8618 ( .A1(n11785), .A2(n7354), .ZN(n14110) );
  NAND2_X1 U8619 ( .A1(n14202), .A2(n11841), .ZN(n14122) );
  NAND2_X1 U8620 ( .A1(n9216), .A2(n9215), .ZN(n14131) );
  NAND2_X1 U8621 ( .A1(n6832), .A2(n11809), .ZN(n6827) );
  AND2_X1 U8622 ( .A1(n14214), .A2(n6830), .ZN(n6829) );
  NAND2_X1 U8623 ( .A1(n6838), .A2(n6837), .ZN(n6836) );
  NAND2_X1 U8624 ( .A1(n6840), .A2(n11885), .ZN(n6839) );
  NAND2_X1 U8625 ( .A1(n14194), .A2(n11831), .ZN(n14148) );
  NAND2_X1 U8626 ( .A1(n14185), .A2(n14184), .ZN(n6655) );
  NAND2_X1 U8627 ( .A1(n14230), .A2(n11795), .ZN(n14167) );
  INV_X1 U8628 ( .A(n14647), .ZN(n14173) );
  INV_X1 U8629 ( .A(n14259), .ZN(n14869) );
  AND4_X1 U8630 ( .A1(n10863), .A2(n10862), .A3(n10861), .A4(n10860), .ZN(
        n11780) );
  AND2_X1 U8631 ( .A1(n14820), .A2(n14821), .ZN(n11022) );
  NAND2_X1 U8632 ( .A1(n8982), .A2(n8981), .ZN(n9211) );
  NAND2_X1 U8633 ( .A1(n6828), .A2(n11809), .ZN(n14213) );
  NAND2_X1 U8634 ( .A1(n14176), .A2(n14177), .ZN(n6828) );
  AND2_X1 U8635 ( .A1(n6854), .A2(n9614), .ZN(n10110) );
  OR2_X1 U8636 ( .A1(n9615), .A2(n7406), .ZN(n6854) );
  AND2_X1 U8637 ( .A1(n9252), .A2(n12178), .ZN(n14883) );
  INV_X1 U8638 ( .A(n14222), .ZN(n6636) );
  AND2_X1 U8639 ( .A1(n14815), .A2(n14961), .ZN(n14879) );
  INV_X1 U8640 ( .A(n14875), .ZN(n14809) );
  OR3_X1 U8641 ( .A1(n11924), .A2(n11923), .A3(n11922), .ZN(n14334) );
  OR2_X1 U8642 ( .A1(n11435), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9000) );
  AND2_X1 U8643 ( .A1(n9081), .A2(n9026), .ZN(n10837) );
  INV_X1 U8644 ( .A(n12159), .ZN(n14552) );
  XNOR2_X1 U8645 ( .A(n11456), .B(n12157), .ZN(n14564) );
  AOI21_X1 U8646 ( .B1(n11763), .B2(n14832), .A(n11762), .ZN(n14569) );
  NAND2_X1 U8647 ( .A1(n11758), .A2(n11759), .ZN(n11763) );
  NAND2_X1 U8648 ( .A1(n6793), .A2(n14832), .ZN(n6626) );
  NAND2_X1 U8649 ( .A1(n14354), .A2(n14729), .ZN(n6792) );
  AND2_X1 U8650 ( .A1(n7249), .A2(n7248), .ZN(n14357) );
  NAND2_X1 U8651 ( .A1(n14431), .A2(n14430), .ZN(n14429) );
  NAND2_X1 U8652 ( .A1(n7255), .A2(n11401), .ZN(n14431) );
  NAND2_X1 U8653 ( .A1(n14458), .A2(n7256), .ZN(n7255) );
  NAND2_X1 U8654 ( .A1(n6778), .A2(n6779), .ZN(n14428) );
  OR2_X1 U8655 ( .A1(n14456), .A2(n14439), .ZN(n6778) );
  NAND2_X1 U8656 ( .A1(n11379), .A2(n11378), .ZN(n14470) );
  NAND2_X1 U8657 ( .A1(n7264), .A2(n7265), .ZN(n14496) );
  AND2_X1 U8658 ( .A1(n11444), .A2(n11443), .ZN(n14515) );
  NAND2_X1 U8659 ( .A1(n7268), .A2(n11352), .ZN(n14512) );
  OR2_X1 U8660 ( .A1(n11351), .A2(n11350), .ZN(n7268) );
  NAND2_X1 U8661 ( .A1(n11180), .A2(n11179), .ZN(n14653) );
  NAND2_X1 U8662 ( .A1(n10833), .A2(n10832), .ZN(n14734) );
  AND2_X1 U8663 ( .A1(n10526), .A2(n10525), .ZN(n10708) );
  NAND2_X1 U8664 ( .A1(n7262), .A2(n10547), .ZN(n10704) );
  NAND2_X1 U8665 ( .A1(n10546), .A2(n10545), .ZN(n7262) );
  INV_X1 U8666 ( .A(n14956), .ZN(n10375) );
  NAND2_X1 U8667 ( .A1(n14544), .A2(n9272), .ZN(n14506) );
  NOR2_X1 U8668 ( .A1(n14743), .A2(n11928), .ZN(n14740) );
  NAND2_X1 U8669 ( .A1(n9685), .A2(n9684), .ZN(n9940) );
  AND2_X1 U8670 ( .A1(n6797), .A2(n6796), .ZN(n6795) );
  NAND2_X1 U8671 ( .A1(n11366), .A2(n9239), .ZN(n6796) );
  NAND2_X1 U8672 ( .A1(n7063), .A2(n6625), .ZN(n6624) );
  AND2_X1 U8673 ( .A1(n9220), .A2(n6522), .ZN(n6864) );
  INV_X1 U8674 ( .A(n9217), .ZN(n6625) );
  NAND2_X1 U8675 ( .A1(n14544), .A2(n9269), .ZN(n14546) );
  OR2_X1 U8676 ( .A1(n14616), .A2(n14615), .ZN(n14669) );
  INV_X1 U8677 ( .A(n14953), .ZN(n14975) );
  NAND2_X1 U8678 ( .A1(n12115), .A2(n12114), .ZN(n14074) );
  INV_X1 U8679 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8689) );
  NAND2_X1 U8680 ( .A1(n7081), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8328) );
  INV_X1 U8681 ( .A(n8163), .ZN(n7076) );
  XNOR2_X1 U8682 ( .A(n11317), .B(n11316), .ZN(n11488) );
  CLKBUF_X1 U8683 ( .A(n14885), .Z(n6663) );
  NAND2_X1 U8684 ( .A1(n8171), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n8176) );
  NOR2_X1 U8685 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n8173) );
  XNOR2_X1 U8686 ( .A(n11403), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14696) );
  INV_X1 U8687 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10087) );
  INV_X1 U8688 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9541) );
  INV_X1 U8689 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9428) );
  INV_X1 U8690 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9083) );
  INV_X1 U8691 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9039) );
  INV_X1 U8692 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n8640) );
  INV_X1 U8693 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8472) );
  INV_X1 U8694 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8377) );
  OAI21_X1 U8695 ( .B1(n8376), .B2(n8375), .A(n8463), .ZN(n10379) );
  INV_X1 U8696 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8365) );
  INV_X1 U8697 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n13735) );
  INV_X1 U8698 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n8308) );
  NOR2_X1 U8699 ( .A1(n15257), .A2(n7485), .ZN(n14706) );
  NAND2_X1 U8700 ( .A1(n14705), .A2(n6751), .ZN(n15254) );
  OAI21_X1 U8701 ( .B1(n14706), .B2(n14707), .A(n6752), .ZN(n6751) );
  INV_X1 U8702 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6752) );
  NOR2_X1 U8703 ( .A1(n15254), .A2(n15255), .ZN(n15253) );
  XNOR2_X1 U8704 ( .A(n7487), .B(n15015), .ZN(n15244) );
  XNOR2_X1 U8705 ( .A(n7490), .B(n6750), .ZN(n15248) );
  NAND2_X1 U8706 ( .A1(n15248), .A2(n15247), .ZN(n15246) );
  NAND2_X1 U8707 ( .A1(n14712), .A2(n7505), .ZN(n7507) );
  OAI21_X1 U8708 ( .B1(n14844), .B2(n14845), .A(n6807), .ZN(n6806) );
  NOR2_X1 U8709 ( .A1(n7516), .A2(n7517), .ZN(n14856) );
  NAND2_X1 U8710 ( .A1(n14860), .A2(n14862), .ZN(n14866) );
  NOR2_X1 U8711 ( .A1(n14866), .A2(n14867), .ZN(n14865) );
  OR2_X1 U8712 ( .A1(n14754), .A2(n6743), .ZN(n6739) );
  INV_X1 U8713 ( .A(n12964), .ZN(n7008) );
  XNOR2_X1 U8714 ( .A(n6587), .B(n6586), .ZN(n13079) );
  INV_X1 U8715 ( .A(n13057), .ZN(n6586) );
  NAND2_X1 U8716 ( .A1(n6706), .A2(n6705), .ZN(P3_U3456) );
  NAND2_X1 U8717 ( .A1(n15234), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n6705) );
  NAND2_X1 U8718 ( .A1(n11670), .A2(n15232), .ZN(n6706) );
  AND2_X1 U8719 ( .A1(n9609), .A2(n9112), .ZN(n9121) );
  OR2_X1 U8720 ( .A1(n7005), .A2(n6611), .ZN(P2_U3236) );
  OAI21_X1 U8721 ( .B1(n13947), .B2(n13871), .A(n6612), .ZN(n6611) );
  OAI21_X1 U8722 ( .B1(n13946), .B2(n15075), .A(n7006), .ZN(n7005) );
  NAND2_X1 U8723 ( .A1(n13943), .A2(n15064), .ZN(n6612) );
  NAND2_X1 U8724 ( .A1(n12177), .A2(n12178), .ZN(n6606) );
  OR2_X1 U8725 ( .A1(n14977), .A2(n7060), .ZN(n7059) );
  NAND2_X1 U8726 ( .A1(n14659), .A2(n14977), .ZN(n7061) );
  INV_X1 U8727 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7060) );
  OAI21_X1 U8728 ( .B1(n14074), .B2(n14694), .A(n7357), .ZN(P1_U3325) );
  NOR2_X1 U8729 ( .A1(n7359), .A2(n7358), .ZN(n7357) );
  NOR2_X1 U8730 ( .A1(n7356), .A2(P1_U3086), .ZN(n7358) );
  NOR2_X1 U8731 ( .A1(n14684), .A2(n12504), .ZN(n7359) );
  NAND2_X1 U8732 ( .A1(n6728), .A2(n6725), .ZN(n15251) );
  INV_X1 U8733 ( .A(n6731), .ZN(n15250) );
  OAI21_X1 U8734 ( .B1(n7497), .B2(n14709), .A(P2_ADDR_REG_7__SCAN_IN), .ZN(
        n6725) );
  INV_X1 U8735 ( .A(n6748), .ZN(n14851) );
  INV_X1 U8736 ( .A(n14862), .ZN(n14861) );
  NAND2_X1 U8737 ( .A1(n6744), .A2(n6740), .ZN(n7532) );
  AND2_X1 U8738 ( .A1(n7188), .A2(n7185), .ZN(n6425) );
  XNOR2_X1 U8739 ( .A(n7525), .B(n7524), .ZN(n14701) );
  INV_X1 U8740 ( .A(n14701), .ZN(n6747) );
  AND2_X1 U8741 ( .A1(n14495), .A2(n7094), .ZN(n6426) );
  AND2_X1 U8742 ( .A1(n7383), .A2(n6442), .ZN(n6427) );
  AND2_X1 U8743 ( .A1(n13305), .A2(n13200), .ZN(n6428) );
  AND2_X1 U8744 ( .A1(n12907), .A2(n7043), .ZN(n6429) );
  AND2_X1 U8745 ( .A1(n7195), .A2(n9912), .ZN(n6430) );
  INV_X1 U8746 ( .A(n13801), .ZN(n7199) );
  NAND2_X1 U8747 ( .A1(n11319), .A2(n11318), .ZN(n14566) );
  OR2_X1 U8748 ( .A1(n12872), .A2(n13163), .ZN(n6431) );
  NAND2_X1 U8749 ( .A1(n11343), .A2(n11342), .ZN(n14403) );
  INV_X1 U8750 ( .A(n14403), .ZN(n6782) );
  AND2_X1 U8751 ( .A1(n7415), .A2(n7599), .ZN(n6432) );
  AND2_X1 U8752 ( .A1(n6787), .A2(n11181), .ZN(n6433) );
  OR2_X1 U8753 ( .A1(n7186), .A2(n13590), .ZN(n6434) );
  NAND2_X1 U8754 ( .A1(n7296), .A2(n7591), .ZN(n7742) );
  AND2_X1 U8755 ( .A1(n8462), .A2(n8288), .ZN(n6435) );
  AND2_X1 U8756 ( .A1(n6785), .A2(n6498), .ZN(n6436) );
  OR2_X1 U8757 ( .A1(n6486), .A2(n7210), .ZN(n6437) );
  OR2_X1 U8758 ( .A1(n7346), .A2(n6942), .ZN(n6438) );
  NAND2_X1 U8759 ( .A1(n11789), .A2(n11790), .ZN(n6439) );
  INV_X1 U8760 ( .A(n7107), .ZN(n7105) );
  AND2_X1 U8761 ( .A1(n7320), .A2(n7319), .ZN(n7107) );
  OR2_X1 U8762 ( .A1(n7893), .A2(n11096), .ZN(n6440) );
  INV_X1 U8763 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8586) );
  NAND4_X1 U8764 ( .A1(n9258), .A2(n9257), .A3(n9256), .A4(n9255), .ZN(n14262)
         );
  AND2_X1 U8765 ( .A1(n7236), .A2(n6491), .ZN(n6441) );
  INV_X1 U8766 ( .A(n13185), .ZN(n13163) );
  AND2_X1 U8767 ( .A1(n12360), .A2(n12359), .ZN(n6442) );
  AND2_X1 U8768 ( .A1(n12241), .A2(n12240), .ZN(n6443) );
  NOR2_X1 U8769 ( .A1(n12314), .A2(n6956), .ZN(n6444) );
  AND2_X1 U8770 ( .A1(n7100), .A2(n7103), .ZN(n6445) );
  INV_X1 U8771 ( .A(n7053), .ZN(n7052) );
  NAND2_X1 U8772 ( .A1(n8056), .A2(n12819), .ZN(n7053) );
  AND2_X1 U8773 ( .A1(n6875), .A2(n6440), .ZN(n13256) );
  INV_X1 U8774 ( .A(n13175), .ZN(n6887) );
  INV_X1 U8775 ( .A(n11692), .ZN(n6764) );
  INV_X1 U8776 ( .A(n12471), .ZN(n7225) );
  INV_X1 U8777 ( .A(n14806), .ZN(n6799) );
  AND2_X1 U8778 ( .A1(n8593), .A2(n14076), .ZN(n6446) );
  INV_X1 U8779 ( .A(n12975), .ZN(n6635) );
  OR2_X1 U8780 ( .A1(n13277), .A2(n12569), .ZN(n12907) );
  AND2_X1 U8781 ( .A1(n7108), .A2(n6445), .ZN(n6447) );
  AND2_X1 U8782 ( .A1(n8491), .A2(n6656), .ZN(n6448) );
  INV_X1 U8783 ( .A(n6446), .ZN(n9352) );
  INV_X1 U8784 ( .A(n9352), .ZN(n10688) );
  INV_X1 U8785 ( .A(n12456), .ZN(n7209) );
  AND2_X1 U8786 ( .A1(n10209), .A2(n10208), .ZN(n6449) );
  AND2_X1 U8787 ( .A1(n12147), .A2(n12024), .ZN(n6450) );
  AND2_X1 U8788 ( .A1(n6999), .A2(n11635), .ZN(n6451) );
  NAND2_X1 U8789 ( .A1(n7609), .A2(n7608), .ZN(n12899) );
  INV_X1 U8790 ( .A(n12460), .ZN(n7197) );
  INV_X1 U8791 ( .A(n9387), .ZN(n11947) );
  INV_X1 U8792 ( .A(n12483), .ZN(n7007) );
  OR2_X1 U8793 ( .A1(n7499), .A2(n7500), .ZN(n6452) );
  AND2_X1 U8794 ( .A1(n12843), .A2(n12837), .ZN(n6453) );
  INV_X1 U8795 ( .A(n6940), .ZN(n6939) );
  INV_X1 U8796 ( .A(n11885), .ZN(n6845) );
  INV_X1 U8797 ( .A(n7163), .ZN(n7162) );
  AND2_X1 U8798 ( .A1(n7307), .A2(n12513), .ZN(n6454) );
  AND2_X1 U8799 ( .A1(n7147), .A2(n6704), .ZN(n6455) );
  AND2_X1 U8800 ( .A1(n7248), .A2(n14373), .ZN(n6457) );
  OR2_X1 U8801 ( .A1(n13780), .A2(n13536), .ZN(n6458) );
  AND2_X1 U8802 ( .A1(n12020), .A2(n12022), .ZN(n12147) );
  NOR2_X1 U8803 ( .A1(n7730), .A2(n7297), .ZN(n7744) );
  NOR2_X1 U8804 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7716) );
  AND2_X1 U8805 ( .A1(n9721), .A2(n9704), .ZN(n6459) );
  INV_X1 U8806 ( .A(n12044), .ZN(n14478) );
  AND2_X1 U8807 ( .A1(n13371), .A2(n12538), .ZN(n6460) );
  OR2_X1 U8808 ( .A1(n13846), .A2(n11694), .ZN(n6461) );
  AND2_X1 U8809 ( .A1(n12907), .A2(n12947), .ZN(n6462) );
  XNOR2_X1 U8810 ( .A(n14572), .B(n11887), .ZN(n14344) );
  INV_X1 U8811 ( .A(n14344), .ZN(n7074) );
  OR2_X1 U8812 ( .A1(n6593), .A2(n13548), .ZN(n6463) );
  OR2_X1 U8813 ( .A1(n14349), .A2(n14243), .ZN(n6464) );
  AND2_X1 U8814 ( .A1(n12308), .A2(n13546), .ZN(n6465) );
  OR2_X1 U8815 ( .A1(n11452), .A2(n14392), .ZN(n6466) );
  INV_X1 U8816 ( .A(n9218), .ZN(n6865) );
  INV_X1 U8817 ( .A(n11977), .ZN(n7124) );
  INV_X1 U8818 ( .A(n12857), .ZN(n7048) );
  OR2_X1 U8819 ( .A1(n12872), .A2(n13185), .ZN(n6467) );
  XOR2_X1 U8820 ( .A(n13064), .B(n13065), .Z(n6468) );
  NAND2_X1 U8821 ( .A1(n7655), .A2(n7415), .ZN(n6469) );
  INV_X1 U8822 ( .A(n12839), .ZN(n7035) );
  OR2_X1 U8823 ( .A1(n11404), .A2(n14274), .ZN(n6470) );
  NAND2_X1 U8824 ( .A1(n12695), .A2(n13175), .ZN(n6471) );
  AND2_X1 U8825 ( .A1(n8166), .A2(n8702), .ZN(n6472) );
  NAND2_X1 U8826 ( .A1(n8591), .A2(n8592), .ZN(n14076) );
  AND2_X1 U8827 ( .A1(n6447), .A2(n12177), .ZN(n6473) );
  AND2_X1 U8828 ( .A1(n7424), .A2(n12171), .ZN(n6474) );
  AND4_X1 U8829 ( .A1(n7640), .A2(n7639), .A3(n7638), .A4(n7637), .ZN(n13175)
         );
  OR2_X1 U8830 ( .A1(n11209), .A2(n11210), .ZN(n6475) );
  AND2_X1 U8831 ( .A1(n12314), .A2(n11230), .ZN(n6476) );
  AND2_X1 U8832 ( .A1(n13954), .A2(n13535), .ZN(n6477) );
  OR2_X1 U8833 ( .A1(n13155), .A2(n13164), .ZN(n12763) );
  INV_X1 U8834 ( .A(n13960), .ZN(n13780) );
  AND2_X1 U8835 ( .A1(n12547), .A2(n13163), .ZN(n6478) );
  NAND2_X1 U8836 ( .A1(n11500), .A2(n11499), .ZN(n13536) );
  AND2_X1 U8837 ( .A1(n12288), .A2(n12287), .ZN(n6479) );
  NAND2_X1 U8838 ( .A1(n11567), .A2(n11566), .ZN(n13973) );
  INV_X1 U8839 ( .A(n12909), .ZN(n13087) );
  AND2_X1 U8840 ( .A1(n12245), .A2(n13554), .ZN(n6480) );
  AND2_X1 U8841 ( .A1(n12332), .A2(n12331), .ZN(n6481) );
  AND2_X1 U8842 ( .A1(n12267), .A2(n12266), .ZN(n6482) );
  INV_X1 U8844 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14068) );
  AND2_X1 U8845 ( .A1(n14606), .A2(n14150), .ZN(n6483) );
  NAND2_X1 U8846 ( .A1(n7206), .A2(n6461), .ZN(n6484) );
  NAND2_X1 U8847 ( .A1(n13601), .A2(n13600), .ZN(n6485) );
  AND2_X1 U8848 ( .A1(n9441), .A2(n7211), .ZN(n6486) );
  INV_X1 U8849 ( .A(n7205), .ZN(n7204) );
  NAND2_X1 U8850 ( .A1(n13827), .A2(n6461), .ZN(n7205) );
  AND2_X1 U8851 ( .A1(n7382), .A2(n7380), .ZN(n6487) );
  AND2_X1 U8852 ( .A1(n12674), .A2(n7301), .ZN(n6488) );
  OR2_X1 U8853 ( .A1(n12228), .A2(n12226), .ZN(n6489) );
  AND2_X1 U8854 ( .A1(n13977), .A2(n13539), .ZN(n6490) );
  NAND2_X1 U8855 ( .A1(n13423), .A2(n13422), .ZN(n6491) );
  AND2_X1 U8856 ( .A1(n14806), .A2(n14257), .ZN(n6492) );
  AND2_X1 U8857 ( .A1(n7225), .A2(n10930), .ZN(n6493) );
  INV_X1 U8858 ( .A(n14331), .ZN(n14555) );
  AND2_X1 U8859 ( .A1(n11450), .A2(n14150), .ZN(n6494) );
  INV_X1 U8860 ( .A(n12873), .ZN(n7020) );
  OR2_X1 U8861 ( .A1(n13305), .A2(n13174), .ZN(n12873) );
  NAND2_X1 U8862 ( .A1(n7104), .A2(n6474), .ZN(n7103) );
  AND2_X1 U8863 ( .A1(n13128), .A2(n13135), .ZN(n6495) );
  AND2_X1 U8864 ( .A1(n11847), .A2(n11846), .ZN(n6496) );
  INV_X1 U8865 ( .A(n11815), .ZN(n6832) );
  INV_X1 U8866 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6657) );
  INV_X1 U8867 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8702) );
  AND2_X1 U8868 ( .A1(n11878), .A2(n11877), .ZN(n6497) );
  OR2_X1 U8869 ( .A1(n7095), .A2(n6786), .ZN(n6498) );
  NOR2_X1 U8870 ( .A1(n14632), .A2(n14638), .ZN(n6499) );
  NOR2_X1 U8871 ( .A1(n14451), .A2(n11448), .ZN(n6500) );
  OR2_X1 U8872 ( .A1(n7383), .A2(n6442), .ZN(n6501) );
  AND4_X1 U8873 ( .A1(n7601), .A2(n8030), .A3(n8069), .A4(n7600), .ZN(n6502)
         );
  AND2_X1 U8874 ( .A1(n7234), .A2(n6441), .ZN(n6503) );
  OR2_X1 U8875 ( .A1(n11642), .A2(n6973), .ZN(n6504) );
  AND2_X1 U8876 ( .A1(n6894), .A2(n8002), .ZN(n6505) );
  NOR2_X1 U8877 ( .A1(n13758), .A2(n7187), .ZN(n7186) );
  INV_X1 U8878 ( .A(n7796), .ZN(n7797) );
  NAND2_X1 U8879 ( .A1(n7716), .A2(n7590), .ZN(n7730) );
  NOR2_X1 U8880 ( .A1(n14636), .A2(n14250), .ZN(n6506) );
  INV_X1 U8881 ( .A(n12039), .ZN(n7095) );
  INV_X1 U8882 ( .A(n12872), .ZN(n13365) );
  NAND2_X1 U8883 ( .A1(n7973), .A2(n7972), .ZN(n12872) );
  AND2_X1 U8884 ( .A1(n12854), .A2(n12853), .ZN(n13237) );
  INV_X1 U8885 ( .A(n8025), .ZN(n6714) );
  AND2_X1 U8886 ( .A1(n12024), .A2(n12023), .ZN(n14534) );
  AND2_X1 U8887 ( .A1(n11869), .A2(n11868), .ZN(n6507) );
  AND2_X1 U8888 ( .A1(n9414), .A2(n9413), .ZN(n6508) );
  AND2_X1 U8889 ( .A1(n8285), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6509) );
  INV_X1 U8890 ( .A(n12695), .ZN(n13361) );
  NAND2_X1 U8891 ( .A1(n7644), .A2(n7643), .ZN(n12695) );
  NAND2_X1 U8892 ( .A1(n12027), .A2(n12026), .ZN(n6510) );
  INV_X1 U8893 ( .A(n6987), .ZN(n6991) );
  OR2_X1 U8894 ( .A1(n10660), .A2(n6992), .ZN(n6987) );
  AND2_X1 U8895 ( .A1(n13361), .A2(n13175), .ZN(n6511) );
  AND2_X1 U8896 ( .A1(n12872), .A2(n13185), .ZN(n6512) );
  AND2_X1 U8897 ( .A1(n12695), .A2(n6887), .ZN(n6513) );
  AND2_X1 U8898 ( .A1(n10187), .A2(n10188), .ZN(n6514) );
  NAND2_X1 U8899 ( .A1(n10925), .A2(n10924), .ZN(n12308) );
  NOR2_X1 U8900 ( .A1(n11862), .A2(n14103), .ZN(n6515) );
  OAI21_X1 U8901 ( .B1(n13188), .B2(n7020), .A(n12877), .ZN(n7019) );
  INV_X1 U8902 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8588) );
  INV_X1 U8903 ( .A(n12242), .ZN(n7390) );
  INV_X1 U8904 ( .A(n12361), .ZN(n7383) );
  NAND2_X1 U8905 ( .A1(n13266), .A2(n7035), .ZN(n6516) );
  NAND2_X1 U8906 ( .A1(n7423), .A2(n6501), .ZN(n6517) );
  AND3_X1 U8907 ( .A1(n8495), .A2(n13732), .A3(n8496), .ZN(n6518) );
  INV_X1 U8908 ( .A(n12314), .ZN(n14065) );
  NAND2_X1 U8909 ( .A1(n11071), .A2(n11070), .ZN(n12314) );
  AND2_X1 U8910 ( .A1(n7100), .A2(n7101), .ZN(n6519) );
  AND2_X1 U8911 ( .A1(n12272), .A2(n12271), .ZN(n6520) );
  OR2_X1 U8912 ( .A1(n12291), .A2(n6479), .ZN(n6521) );
  OR2_X1 U8913 ( .A1(n11404), .A2(n6865), .ZN(n6522) );
  OR2_X1 U8914 ( .A1(n6842), .A2(n6845), .ZN(n6523) );
  AND2_X1 U8915 ( .A1(n7505), .A2(n6737), .ZN(n6524) );
  NOR2_X1 U8916 ( .A1(n14835), .A2(n14254), .ZN(n6525) );
  NOR2_X1 U8917 ( .A1(n7319), .A2(n7320), .ZN(n6526) );
  INV_X1 U8918 ( .A(n6893), .ZN(n6892) );
  NOR2_X1 U8919 ( .A1(n12926), .A2(n6724), .ZN(n6893) );
  NAND2_X1 U8920 ( .A1(n7655), .A2(n7310), .ZN(n6527) );
  NOR2_X1 U8921 ( .A1(n13140), .A2(n12764), .ZN(n6528) );
  AND2_X1 U8922 ( .A1(n7382), .A2(n12357), .ZN(n6529) );
  AND2_X1 U8923 ( .A1(n11181), .A2(n11176), .ZN(n6530) );
  OR2_X1 U8924 ( .A1(n12057), .A2(n12055), .ZN(n6531) );
  INV_X1 U8925 ( .A(n6906), .ZN(n6905) );
  NAND2_X1 U8926 ( .A1(n13239), .A2(n13221), .ZN(n6906) );
  OR2_X1 U8927 ( .A1(n7392), .A2(n6481), .ZN(n6532) );
  AND2_X1 U8928 ( .A1(n7374), .A2(n8691), .ZN(n6533) );
  NAND2_X1 U8929 ( .A1(n12086), .A2(n7122), .ZN(n6534) );
  INV_X1 U8930 ( .A(n7189), .ZN(n7188) );
  NAND2_X1 U8931 ( .A1(n6458), .A2(n7190), .ZN(n7189) );
  NAND2_X1 U8932 ( .A1(n11997), .A2(n7119), .ZN(n6535) );
  INV_X1 U8933 ( .A(n11642), .ZN(n6975) );
  INV_X1 U8934 ( .A(n7417), .ZN(n6873) );
  OR2_X1 U8935 ( .A1(n7390), .A2(n6443), .ZN(n6536) );
  OR2_X1 U8936 ( .A1(n12311), .A2(n6541), .ZN(n6537) );
  INV_X1 U8937 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8327) );
  INV_X1 U8938 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n8204) );
  INV_X1 U8939 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n13734) );
  INV_X1 U8940 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6771) );
  INV_X1 U8941 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8495) );
  AND3_X1 U8942 ( .A1(n6607), .A2(n6606), .A3(n7098), .ZN(P1_U3242) );
  INV_X1 U8943 ( .A(n13459), .ZN(n13424) );
  INV_X1 U8944 ( .A(n9173), .ZN(n6583) );
  NAND2_X1 U8945 ( .A1(n11095), .A2(n7894), .ZN(n6875) );
  INV_X1 U8946 ( .A(n6924), .ZN(n6923) );
  NAND2_X1 U8947 ( .A1(n11159), .A2(n6925), .ZN(n6924) );
  XOR2_X1 U8948 ( .A(n11876), .B(n11877), .Z(n6539) );
  AOI21_X1 U8949 ( .B1(n13232), .B2(n13231), .A(n6905), .ZN(n13220) );
  XOR2_X1 U8950 ( .A(n11794), .B(n11793), .Z(n6540) );
  NAND2_X1 U8951 ( .A1(n10596), .A2(n8051), .ZN(n10811) );
  OR2_X1 U8952 ( .A1(n14017), .A2(n10562), .ZN(n10662) );
  INV_X1 U8953 ( .A(n10662), .ZN(n6955) );
  INV_X1 U8954 ( .A(n14345), .ZN(n12097) );
  NAND2_X1 U8955 ( .A1(n10526), .A2(n7093), .ZN(n10707) );
  NAND2_X1 U8956 ( .A1(n11444), .A2(n7096), .ZN(n14513) );
  NAND4_X1 U8957 ( .A1(n11324), .A2(n11323), .A3(n11322), .A4(n11321), .ZN(
        n14243) );
  AND2_X1 U8958 ( .A1(n12307), .A2(n12306), .ZN(n6541) );
  AND2_X1 U8959 ( .A1(n12566), .A2(n12565), .ZN(n6542) );
  AND2_X1 U8960 ( .A1(n10559), .A2(n10558), .ZN(n6543) );
  INV_X1 U8961 ( .A(n6949), .ZN(n13897) );
  NOR2_X1 U8962 ( .A1(n13898), .A2(n13899), .ZN(n6949) );
  AND2_X1 U8963 ( .A1(n6789), .A2(n12024), .ZN(n6544) );
  INV_X1 U8964 ( .A(n11330), .ZN(n7342) );
  AND2_X1 U8965 ( .A1(n6900), .A2(n6899), .ZN(n6545) );
  INV_X1 U8966 ( .A(n11809), .ZN(n6831) );
  OR2_X1 U8967 ( .A1(n11808), .A2(n11807), .ZN(n11809) );
  AND2_X1 U8968 ( .A1(n7000), .A2(n6451), .ZN(n6546) );
  AND2_X1 U8969 ( .A1(n10359), .A2(n10358), .ZN(n6547) );
  AND2_X1 U8970 ( .A1(n12341), .A2(n12340), .ZN(n6548) );
  INV_X1 U8971 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7610) );
  AND2_X1 U8972 ( .A1(n7036), .A2(n7035), .ZN(n6549) );
  AND2_X1 U8973 ( .A1(n10880), .A2(n12819), .ZN(n6550) );
  OR2_X1 U8974 ( .A1(n12344), .A2(n6548), .ZN(n6551) );
  INV_X1 U8975 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9045) );
  AND2_X1 U8976 ( .A1(n8126), .A2(n8125), .ZN(n15234) );
  NAND2_X1 U8977 ( .A1(n11514), .A2(n11513), .ZN(n13881) );
  INV_X1 U8978 ( .A(n13881), .ZN(n6948) );
  INV_X1 U8979 ( .A(n12294), .ZN(n6959) );
  INV_X1 U8980 ( .A(n7339), .ZN(n7337) );
  NOR2_X1 U8981 ( .A1(n11424), .A2(n7340), .ZN(n7339) );
  AND2_X1 U8982 ( .A1(n9482), .A2(n9481), .ZN(n6552) );
  AND2_X1 U8983 ( .A1(n7276), .A2(n7274), .ZN(n6553) );
  AND2_X1 U8984 ( .A1(n11538), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U8985 ( .A1(n9593), .A2(n6420), .ZN(n6555) );
  AND2_X1 U8986 ( .A1(n11292), .A2(n12511), .ZN(n6556) );
  AND2_X1 U8987 ( .A1(n7574), .A2(n11512), .ZN(n6557) );
  INV_X1 U8988 ( .A(n13262), .ZN(n6878) );
  NAND2_X1 U8989 ( .A1(n8786), .A2(n8785), .ZN(n14832) );
  INV_X1 U8990 ( .A(n11973), .ZN(n7091) );
  XNOR2_X1 U8991 ( .A(n7946), .B(n7945), .ZN(n13044) );
  INV_X1 U8992 ( .A(n15093), .ZN(n14012) );
  INV_X1 U8993 ( .A(n12268), .ZN(n6950) );
  INV_X1 U8994 ( .A(SI_24_), .ZN(n6925) );
  INV_X1 U8995 ( .A(n8045), .ZN(n13056) );
  NAND2_X1 U8996 ( .A1(n9624), .A2(n9623), .ZN(n6558) );
  INV_X1 U8997 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11565) );
  AND2_X1 U8998 ( .A1(n14081), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6559) );
  INV_X1 U8999 ( .A(n7228), .ZN(n9725) );
  NOR2_X1 U9000 ( .A1(n11651), .A2(n7176), .ZN(n7175) );
  INV_X1 U9001 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n6807) );
  AND2_X1 U9002 ( .A1(n12440), .A2(n12439), .ZN(n6560) );
  INV_X1 U9003 ( .A(n13044), .ZN(n6581) );
  NAND2_X1 U9004 ( .A1(n9929), .A2(n9944), .ZN(n10270) );
  NAND2_X1 U9005 ( .A1(n10378), .A2(n10377), .ZN(n10546) );
  NAND2_X1 U9006 ( .A1(n9390), .A2(n7420), .ZN(n9517) );
  NAND2_X1 U9007 ( .A1(n7421), .A2(n10972), .ZN(n11177) );
  OAI22_X1 U9008 ( .A1(n14477), .A2(n12044), .B1(n14248), .B2(n14489), .ZN(
        n14460) );
  OAI22_X1 U9009 ( .A1(n9922), .A2(n12134), .B1(n14262), .B2(n11973), .ZN(
        n10005) );
  NAND2_X1 U9010 ( .A1(n11351), .A2(n7266), .ZN(n7264) );
  NAND2_X1 U9011 ( .A1(n14411), .A2(n14410), .ZN(n14409) );
  NAND3_X2 U9012 ( .A1(n8790), .A2(n6561), .A3(n8792), .ZN(n14265) );
  NOR2_X1 U9013 ( .A1(n14342), .A2(n6944), .ZN(n11765) );
  NAND3_X2 U9014 ( .A1(n8700), .A2(n6562), .A3(n8699), .ZN(n14267) );
  AND2_X1 U9015 ( .A1(n8701), .A2(n8698), .ZN(n6562) );
  AND2_X2 U9016 ( .A1(n7356), .A2(n8693), .ZN(n8996) );
  XNOR2_X2 U9017 ( .A(n8690), .B(n8689), .ZN(n7356) );
  NAND2_X1 U9018 ( .A1(n9394), .A2(n9393), .ZN(n9680) );
  OAI21_X1 U9019 ( .B1(n14403), .B2(n14244), .A(n14391), .ZN(n14372) );
  OAI22_X1 U9020 ( .A1(n10829), .A2(n10828), .B1(n14256), .B2(n14828), .ZN(
        n14721) );
  MUX2_X1 U9021 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14659), .S(n14986), .Z(
        P1_U3557) );
  NAND2_X1 U9022 ( .A1(n9517), .A2(n9516), .ZN(n9392) );
  OAI21_X2 U9023 ( .B1(n8325), .B2(n7376), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8692) );
  NAND2_X2 U9024 ( .A1(n11715), .A2(n10717), .ZN(n11063) );
  NAND2_X1 U9025 ( .A1(n8468), .A2(n8632), .ZN(n10527) );
  NAND2_X1 U9026 ( .A1(n10078), .A2(n10077), .ZN(n6563) );
  NAND2_X1 U9027 ( .A1(n6426), .A2(n6785), .ZN(n6784) );
  OAI21_X2 U9028 ( .B1(n9697), .B2(n7242), .A(n7240), .ZN(n9848) );
  NAND2_X1 U9029 ( .A1(n6602), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7425) );
  NAND2_X1 U9030 ( .A1(n11704), .A2(n6759), .ZN(n11715) );
  NOR2_X1 U9031 ( .A1(n14848), .A2(n14849), .ZN(n14847) );
  NAND2_X1 U9032 ( .A1(n6748), .A2(n6576), .ZN(n7516) );
  NAND2_X1 U9033 ( .A1(n14853), .A2(n14852), .ZN(n6749) );
  AND2_X2 U9034 ( .A1(n14855), .A2(n14857), .ZN(n7519) );
  INV_X1 U9035 ( .A(n7491), .ZN(n6750) );
  NAND2_X1 U9036 ( .A1(n14843), .A2(n6806), .ZN(n14848) );
  NAND2_X1 U9037 ( .A1(n14752), .A2(n7523), .ZN(n14700) );
  AOI21_X1 U9038 ( .B1(n7511), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n14847), .ZN(
        n14853) );
  INV_X1 U9039 ( .A(n12297), .ZN(n6567) );
  NAND2_X1 U9040 ( .A1(n12226), .A2(n12228), .ZN(n7398) );
  NAND3_X1 U9041 ( .A1(n6568), .A2(n7379), .A3(n7381), .ZN(n6666) );
  NAND2_X1 U9042 ( .A1(n12358), .A2(n6529), .ZN(n6568) );
  INV_X1 U9043 ( .A(n12222), .ZN(n6596) );
  XNOR2_X1 U9044 ( .A(n6569), .B(n14540), .ZN(n12169) );
  NAND4_X1 U9045 ( .A1(n12158), .A2(n7424), .A3(n12156), .A4(n12157), .ZN(
        n6569) );
  INV_X1 U9046 ( .A(n12172), .ZN(n7108) );
  NAND2_X1 U9047 ( .A1(n6599), .A2(n6915), .ZN(n11288) );
  NAND2_X1 U9048 ( .A1(n7341), .A2(n7338), .ZN(n11425) );
  NAND2_X1 U9049 ( .A1(n9587), .A2(n9586), .ZN(n10078) );
  NAND2_X1 U9050 ( .A1(n7028), .A2(n7027), .ZN(n13236) );
  INV_X1 U9051 ( .A(n7040), .ZN(n12741) );
  INV_X1 U9052 ( .A(n7049), .ZN(n13196) );
  NAND2_X1 U9053 ( .A1(n7308), .A2(n7057), .ZN(n7603) );
  NAND2_X1 U9054 ( .A1(n7023), .A2(n7021), .ZN(n10995) );
  NAND2_X1 U9055 ( .A1(n6710), .A2(n6707), .ZN(n11670) );
  OAI21_X1 U9056 ( .B1(n8055), .B2(n7053), .A(n7050), .ZN(n11093) );
  AOI21_X1 U9057 ( .B1(n7056), .B2(n7055), .A(n8061), .ZN(n13107) );
  NAND2_X1 U9058 ( .A1(n6570), .A2(n7139), .ZN(n7138) );
  NAND2_X1 U9059 ( .A1(n12037), .A2(n12036), .ZN(n6570) );
  INV_X1 U9060 ( .A(n7145), .ZN(n12019) );
  NAND2_X1 U9061 ( .A1(n7114), .A2(n7113), .ZN(n12104) );
  NAND2_X1 U9062 ( .A1(n12075), .A2(n12074), .ZN(n12079) );
  NAND2_X1 U9063 ( .A1(n12048), .A2(n12047), .ZN(n12052) );
  NAND2_X1 U9064 ( .A1(n6935), .A2(n6936), .ZN(n6571) );
  INV_X1 U9065 ( .A(n9027), .ZN(n7345) );
  OAI21_X1 U9066 ( .B1(n7346), .B2(n6941), .A(n7344), .ZN(n6940) );
  NAND2_X2 U9067 ( .A1(n10270), .A2(n10269), .ZN(n10376) );
  NAND2_X1 U9068 ( .A1(n11764), .A2(n6622), .ZN(n6621) );
  OAI21_X1 U9069 ( .B1(n9680), .B2(n9679), .A(n9681), .ZN(n9922) );
  NAND2_X1 U9070 ( .A1(n6574), .A2(n6573), .ZN(n6632) );
  NAND2_X1 U9071 ( .A1(n12297), .A2(n12296), .ZN(n6574) );
  INV_X1 U9072 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n8157) );
  INV_X1 U9073 ( .A(n11952), .ZN(n9388) );
  NAND2_X1 U9074 ( .A1(n11183), .A2(n11182), .ZN(n11351) );
  NAND2_X1 U9075 ( .A1(n14858), .A2(n14859), .ZN(n14855) );
  NAND2_X1 U9076 ( .A1(n6749), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6576) );
  NAND2_X1 U9077 ( .A1(n14863), .A2(n14864), .ZN(n14860) );
  NOR2_X1 U9078 ( .A1(n15245), .A2(n15244), .ZN(n15243) );
  NAND2_X1 U9079 ( .A1(n6578), .A2(n6577), .ZN(n6727) );
  INV_X1 U9080 ( .A(n15252), .ZN(n6577) );
  NAND2_X1 U9081 ( .A1(n7497), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6578) );
  NAND2_X1 U9082 ( .A1(n7516), .A2(n7517), .ZN(n14858) );
  NAND4_X1 U9083 ( .A1(n7315), .A2(n7316), .A3(n7314), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7313) );
  NAND2_X1 U9084 ( .A1(n7476), .A2(n8721), .ZN(n6819) );
  INV_X1 U9085 ( .A(n7519), .ZN(n6733) );
  OAI22_X1 U9086 ( .A1(n9367), .A2(n9366), .B1(n9365), .B2(n9375), .ZN(n9976)
         );
  OAI21_X1 U9087 ( .B1(n10154), .B2(n15149), .A(n15143), .ZN(n10335) );
  NAND2_X1 U9088 ( .A1(n13055), .A2(n13058), .ZN(n6588) );
  INV_X1 U9089 ( .A(n13054), .ZN(n6589) );
  NAND2_X1 U9090 ( .A1(n14995), .A2(n8615), .ZN(n6591) );
  NAND2_X1 U9091 ( .A1(n6592), .A2(n10464), .ZN(n10629) );
  NAND2_X1 U9092 ( .A1(n10463), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6592) );
  INV_X4 U9093 ( .A(n13056), .ZN(n13037) );
  NOR2_X1 U9094 ( .A1(n13012), .A2(n13011), .ZN(n13028) );
  NAND2_X1 U9095 ( .A1(n6596), .A2(n6595), .ZN(n6594) );
  NAND2_X1 U9096 ( .A1(n7282), .A2(n7280), .ZN(n12650) );
  NAND2_X1 U9097 ( .A1(n10611), .A2(n10610), .ZN(n7295) );
  NAND2_X1 U9098 ( .A1(n10731), .A2(n10730), .ZN(n10734) );
  NAND2_X1 U9099 ( .A1(n10954), .A2(n10953), .ZN(n10958) );
  OAI21_X1 U9100 ( .B1(n12683), .B2(n12524), .A(n12523), .ZN(n12574) );
  OAI21_X1 U9101 ( .B1(n12531), .B2(n12530), .A(n12529), .ZN(n12658) );
  OAI21_X2 U9102 ( .B1(n7271), .B2(n10058), .A(n7269), .ZN(n10090) );
  NAND2_X1 U9103 ( .A1(n10617), .A2(n10728), .ZN(n10731) );
  NAND2_X1 U9104 ( .A1(n6603), .A2(n6768), .ZN(n10410) );
  NAND2_X1 U9105 ( .A1(n6857), .A2(n6439), .ZN(n7353) );
  NOR2_X1 U9106 ( .A1(n9242), .A2(n9241), .ZN(n9301) );
  NAND2_X1 U9107 ( .A1(n12270), .A2(n7395), .ZN(n7393) );
  NAND2_X1 U9108 ( .A1(n12264), .A2(n12265), .ZN(n12270) );
  NAND3_X1 U9109 ( .A1(n6670), .A2(n7398), .A3(n6594), .ZN(n6628) );
  NAND2_X1 U9110 ( .A1(n6598), .A2(n11944), .ZN(n11951) );
  NAND2_X1 U9111 ( .A1(n11940), .A2(n11941), .ZN(n6598) );
  OAI22_X2 U9112 ( .A1(n7129), .A2(n6456), .B1(n11987), .B2(n7131), .ZN(n11990) );
  OAI22_X2 U9113 ( .A1(n12067), .A2(n7133), .B1(n12066), .B2(n7132), .ZN(
        n12070) );
  NAND2_X2 U9114 ( .A1(n8762), .A2(n8763), .ZN(n14540) );
  INV_X1 U9115 ( .A(n7112), .ZN(n7111) );
  INV_X1 U9116 ( .A(n8167), .ZN(n8760) );
  NAND2_X1 U9117 ( .A1(n8207), .A2(n8266), .ZN(n8231) );
  NAND2_X1 U9118 ( .A1(n10090), .A2(n10091), .ZN(n10262) );
  INV_X1 U9119 ( .A(n9853), .ZN(n9856) );
  INV_X1 U9120 ( .A(n8174), .ZN(n8177) );
  NAND2_X1 U9121 ( .A1(n14157), .A2(n14158), .ZN(n7361) );
  AOI21_X1 U9122 ( .B1(n11005), .B2(n11004), .A(n11003), .ZN(n11008) );
  NAND2_X1 U9123 ( .A1(n7361), .A2(n11861), .ZN(n6637) );
  NAND2_X1 U9124 ( .A1(n8167), .A2(n6472), .ZN(n8322) );
  OAI21_X1 U9125 ( .B1(n12032), .B2(n12031), .A(n12029), .ZN(n12030) );
  NAND2_X1 U9126 ( .A1(n6614), .A2(n7117), .ZN(n12000) );
  NAND2_X1 U9127 ( .A1(n11943), .A2(n7420), .ZN(n11944) );
  NAND2_X1 U9128 ( .A1(n7127), .A2(n7126), .ZN(n11981) );
  OAI21_X1 U9129 ( .B1(n12052), .B2(n12051), .A(n12050), .ZN(n12054) );
  XNOR2_X2 U9130 ( .A(n7522), .B(n6809), .ZN(n14754) );
  NAND2_X1 U9131 ( .A1(n6739), .A2(n6738), .ZN(n14699) );
  XNOR2_X1 U9132 ( .A(n11008), .B(n11010), .ZN(n14873) );
  NAND2_X1 U9133 ( .A1(n7479), .A2(n7478), .ZN(n6815) );
  INV_X1 U9134 ( .A(n7523), .ZN(n6743) );
  AOI21_X1 U9135 ( .B1(n14709), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6727), .ZN(
        n6726) );
  INV_X1 U9136 ( .A(n14865), .ZN(n6811) );
  NAND2_X1 U9137 ( .A1(n6929), .A2(n6927), .ZN(n10744) );
  NAND2_X1 U9138 ( .A1(n6519), .A2(n12177), .ZN(n7099) );
  NAND2_X1 U9139 ( .A1(n11294), .A2(n11293), .ZN(n11317) );
  INV_X1 U9140 ( .A(n7103), .ZN(n7102) );
  NAND2_X1 U9141 ( .A1(n7105), .A2(n6526), .ZN(n7104) );
  INV_X1 U9142 ( .A(n12126), .ZN(n7320) );
  NAND2_X1 U9143 ( .A1(n7229), .A2(n9856), .ZN(n6603) );
  NAND3_X1 U9144 ( .A1(n8366), .A2(n8368), .A3(n8157), .ZN(n8635) );
  INV_X2 U9145 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U9146 ( .A1(n9211), .A2(n9210), .ZN(n9216) );
  NAND2_X1 U9147 ( .A1(n8712), .A2(n8713), .ZN(n8715) );
  NAND2_X1 U9148 ( .A1(n8305), .A2(n8350), .ZN(n9925) );
  OAI21_X1 U9149 ( .B1(n8236), .B2(P2_DATAO_REG_2__SCAN_IN), .A(n6605), .ZN(
        n8220) );
  XNOR2_X1 U9150 ( .A(n6637), .B(n6636), .ZN(n14229) );
  OAI21_X2 U9151 ( .B1(n9301), .B2(n9300), .A(n9299), .ZN(n9615) );
  OR3_X2 U9152 ( .A1(n7321), .A2(n12172), .A3(n7099), .ZN(n6607) );
  NAND2_X2 U9153 ( .A1(n10971), .A2(n10970), .ZN(n14119) );
  NAND2_X1 U9154 ( .A1(n6608), .A2(n9780), .ZN(n9784) );
  XNOR2_X1 U9155 ( .A(n10055), .B(n9779), .ZN(n6608) );
  NAND2_X1 U9156 ( .A1(n12190), .A2(n12189), .ZN(n12197) );
  NOR2_X2 U9157 ( .A1(n9819), .A2(n9785), .ZN(n10058) );
  NAND2_X1 U9158 ( .A1(n7219), .A2(n7218), .ZN(n13858) );
  NAND2_X1 U9159 ( .A1(n6841), .A2(n7360), .ZN(n6650) );
  XNOR2_X1 U9160 ( .A(n6650), .B(n6539), .ZN(n14108) );
  NAND3_X2 U9161 ( .A1(n6654), .A2(n14692), .A3(n8347), .ZN(n9248) );
  NAND2_X1 U9162 ( .A1(n6692), .A2(n12350), .ZN(n12354) );
  NAND3_X1 U9163 ( .A1(n8597), .A2(n6615), .A3(n8594), .ZN(n12180) );
  OAI21_X2 U9164 ( .B1(n7969), .B2(n7180), .A(n7178), .ZN(n7983) );
  NAND2_X1 U9165 ( .A1(n7885), .A2(n7559), .ZN(n7560) );
  NAND2_X2 U9166 ( .A1(n7543), .A2(n7542), .ZN(n7762) );
  NAND2_X1 U9167 ( .A1(n9609), .A2(n7232), .ZN(n9329) );
  OAI21_X1 U9168 ( .B1(n7583), .B2(n7171), .A(n7586), .ZN(n7170) );
  NAND2_X1 U9169 ( .A1(n6955), .A2(n6444), .ZN(n11242) );
  NAND2_X1 U9170 ( .A1(n6949), .A2(n6948), .ZN(n13879) );
  NAND2_X1 U9171 ( .A1(n7308), .A2(n7655), .ZN(n6913) );
  NAND2_X1 U9172 ( .A1(n13842), .A2(n14047), .ZN(n13843) );
  NAND2_X1 U9173 ( .A1(n10367), .A2(n10363), .ZN(n10562) );
  AND2_X2 U9174 ( .A1(n10318), .A2(n15068), .ZN(n9498) );
  NOR2_X2 U9175 ( .A1(n13775), .A2(n13954), .ZN(n11628) );
  NAND3_X1 U9176 ( .A1(n11995), .A2(n6535), .A3(n11994), .ZN(n6614) );
  NAND2_X1 U9177 ( .A1(n8631), .A2(n7324), .ZN(n8632) );
  NAND2_X1 U9178 ( .A1(n7121), .A2(n7120), .ZN(n12090) );
  NAND2_X1 U9179 ( .A1(n6775), .A2(n6774), .ZN(n14415) );
  NAND2_X1 U9180 ( .A1(n12211), .A2(n12210), .ZN(n12217) );
  AOI21_X2 U9181 ( .B1(n12438), .B2(n12437), .A(n12436), .ZN(n12490) );
  NAND2_X1 U9182 ( .A1(n12252), .A2(n12251), .ZN(n12258) );
  AOI21_X1 U9183 ( .B1(n12339), .B2(n12338), .A(n12336), .ZN(n12337) );
  NAND2_X1 U9184 ( .A1(n6619), .A2(n6618), .ZN(n12350) );
  NAND2_X1 U9185 ( .A1(n6617), .A2(n6616), .ZN(n12285) );
  NAND2_X1 U9186 ( .A1(n7399), .A2(n7400), .ZN(n12349) );
  INV_X1 U9187 ( .A(n12349), .ZN(n6619) );
  NAND2_X1 U9188 ( .A1(n9502), .A2(n9504), .ZN(n9394) );
  NOR2_X1 U9189 ( .A1(n6665), .A2(n6664), .ZN(n14342) );
  NAND2_X2 U9190 ( .A1(n14683), .A2(n14885), .ZN(n11404) );
  NAND3_X1 U9191 ( .A1(n7078), .A2(n7076), .A3(n7077), .ZN(n7081) );
  NAND2_X1 U9192 ( .A1(n7244), .A2(n7245), .ZN(n14343) );
  AOI21_X1 U9193 ( .B1(n10967), .B2(n12144), .A(n6525), .ZN(n7421) );
  NAND2_X1 U9194 ( .A1(n6623), .A2(n6533), .ZN(n14677) );
  INV_X1 U9195 ( .A(n8325), .ZN(n6623) );
  OAI21_X1 U9196 ( .B1(n13473), .B2(n11692), .A(n6681), .ZN(n6680) );
  NAND2_X1 U9197 ( .A1(n9329), .A2(n9328), .ZN(n9881) );
  NAND2_X1 U9198 ( .A1(n9592), .A2(n8140), .ZN(n8575) );
  BUF_X1 U9199 ( .A(n13459), .Z(n6627) );
  NAND2_X1 U9200 ( .A1(n6628), .A2(n6489), .ZN(n12234) );
  NAND2_X1 U9201 ( .A1(n12180), .A2(n12432), .ZN(n12184) );
  NAND2_X1 U9202 ( .A1(n6632), .A2(n6631), .ZN(n12303) );
  AOI21_X1 U9203 ( .B1(n12303), .B2(n12302), .A(n12301), .ZN(n12305) );
  NAND3_X1 U9204 ( .A1(n7387), .A2(n6537), .A3(n7386), .ZN(n6639) );
  INV_X1 U9205 ( .A(n12339), .ZN(n6634) );
  NAND2_X1 U9206 ( .A1(n6679), .A2(n7391), .ZN(n12339) );
  NAND2_X1 U9207 ( .A1(n7388), .A2(n7389), .ZN(n12250) );
  XNOR2_X2 U9208 ( .A(n8590), .B(n8589), .ZN(n14073) );
  NAND2_X1 U9209 ( .A1(n7594), .A2(n7773), .ZN(n7878) );
  NAND2_X1 U9210 ( .A1(n12574), .A2(n7284), .ZN(n7282) );
  NOR2_X1 U9211 ( .A1(n8174), .A2(n8173), .ZN(n8175) );
  NAND2_X1 U9212 ( .A1(n6686), .A2(n12419), .ZN(n12438) );
  NAND2_X1 U9213 ( .A1(n6639), .A2(n7385), .ZN(n12318) );
  NAND2_X1 U9214 ( .A1(n12319), .A2(n7403), .ZN(n12325) );
  NAND2_X1 U9215 ( .A1(n8621), .A2(n8478), .ZN(n15004) );
  NAND3_X1 U9216 ( .A1(n12286), .A2(n12285), .A3(n6521), .ZN(n6653) );
  INV_X1 U9217 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n13632) );
  NAND2_X1 U9218 ( .A1(n6646), .A2(n6643), .ZN(n13576) );
  NAND2_X1 U9219 ( .A1(n6644), .A2(n13603), .ZN(n6643) );
  OAI21_X1 U9220 ( .B1(n13571), .B2(n15046), .A(n6645), .ZN(n6644) );
  NAND2_X1 U9221 ( .A1(n13575), .A2(n13574), .ZN(n6646) );
  NAND2_X1 U9222 ( .A1(n9848), .A2(n9847), .ZN(n9853) );
  NOR2_X2 U9223 ( .A1(n11719), .A2(n11718), .ZN(n11723) );
  INV_X1 U9224 ( .A(n7243), .ZN(n7242) );
  AND2_X1 U9225 ( .A1(n11745), .A2(n10206), .ZN(n10207) );
  INV_X1 U9226 ( .A(n14556), .ZN(n14562) );
  NAND2_X1 U9227 ( .A1(n14745), .A2(n14737), .ZN(n14735) );
  NAND2_X1 U9228 ( .A1(n7061), .A2(n7059), .ZN(P1_U3525) );
  INV_X1 U9229 ( .A(n6801), .ZN(n14462) );
  AND2_X2 U9230 ( .A1(n14465), .A2(n14614), .ZN(n14447) );
  OR2_X1 U9231 ( .A1(n10008), .A2(n14944), .ZN(n10009) );
  NOR2_X2 U9232 ( .A1(n14119), .A2(n10976), .ZN(n14531) );
  NOR2_X2 U9233 ( .A1(n14361), .A2(n14572), .ZN(n14348) );
  NAND2_X1 U9234 ( .A1(n6652), .A2(n7128), .ZN(n12062) );
  NAND3_X1 U9235 ( .A1(n12054), .A2(n12053), .A3(n6531), .ZN(n6652) );
  NAND2_X1 U9236 ( .A1(n7138), .A2(n7136), .ZN(n12048) );
  INV_X1 U9237 ( .A(n12104), .ZN(n12107) );
  XNOR2_X2 U9238 ( .A(n9079), .B(n9078), .ZN(n10968) );
  NAND2_X1 U9239 ( .A1(n7323), .A2(n7322), .ZN(n7321) );
  NAND2_X1 U9240 ( .A1(n12070), .A2(n12071), .ZN(n12069) );
  NAND2_X1 U9241 ( .A1(n6653), .A2(n7401), .ZN(n12297) );
  INV_X1 U9242 ( .A(n11164), .ZN(n6654) );
  AND2_X2 U9243 ( .A1(n8181), .A2(n9422), .ZN(n8167) );
  NAND2_X2 U9244 ( .A1(n6655), .A2(n11854), .ZN(n14157) );
  NAND2_X1 U9245 ( .A1(n6849), .A2(n6847), .ZN(n14092) );
  XNOR2_X1 U9246 ( .A(n13001), .B(n11272), .ZN(n11273) );
  NAND2_X2 U9247 ( .A1(n13788), .A2(n11589), .ZN(n13772) );
  NAND2_X1 U9248 ( .A1(n13946), .A2(n6658), .ZN(n14029) );
  NAND2_X2 U9249 ( .A1(n13858), .A2(n11536), .ZN(n13835) );
  NAND2_X1 U9250 ( .A1(n7194), .A2(n7193), .ZN(n10245) );
  XNOR2_X1 U9251 ( .A(n12259), .B(n13553), .ZN(n12460) );
  NAND2_X1 U9252 ( .A1(n8234), .A2(n8233), .ZN(n7318) );
  INV_X1 U9253 ( .A(n10416), .ZN(n6683) );
  NAND2_X1 U9254 ( .A1(n12199), .A2(n12198), .ZN(n12206) );
  INV_X1 U9255 ( .A(n12337), .ZN(n6668) );
  OAI21_X2 U9256 ( .B1(n10376), .B2(n10375), .A(n14869), .ZN(n10378) );
  NAND2_X1 U9257 ( .A1(n6666), .A2(n6687), .ZN(n6686) );
  NAND3_X1 U9258 ( .A1(n6668), .A2(n6669), .A3(n6551), .ZN(n7399) );
  NAND2_X1 U9259 ( .A1(n12258), .A2(n12257), .ZN(n12263) );
  NAND2_X1 U9260 ( .A1(n12222), .A2(n12221), .ZN(n6672) );
  NAND2_X1 U9261 ( .A1(n6672), .A2(n6671), .ZN(n6670) );
  NAND2_X1 U9262 ( .A1(n6678), .A2(n6677), .ZN(n6698) );
  INV_X1 U9263 ( .A(n12318), .ZN(n6674) );
  NAND2_X1 U9264 ( .A1(n6676), .A2(n6675), .ZN(n12286) );
  NAND2_X1 U9265 ( .A1(n12284), .A2(n12283), .ZN(n6676) );
  NAND2_X1 U9266 ( .A1(n12325), .A2(n12326), .ZN(n12324) );
  NAND3_X1 U9267 ( .A1(n12330), .A2(n12329), .A3(n6532), .ZN(n6679) );
  INV_X1 U9268 ( .A(n12215), .ZN(n6696) );
  INV_X1 U9269 ( .A(n6680), .ZN(n11717) );
  INV_X1 U9270 ( .A(n11693), .ZN(n6681) );
  NAND2_X1 U9271 ( .A1(n6760), .A2(n13489), .ZN(n13473) );
  INV_X2 U9272 ( .A(n8236), .ZN(n8968) );
  MUX2_X1 U9273 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8236), .Z(n6943) );
  INV_X1 U9274 ( .A(n8243), .ZN(n8241) );
  NAND2_X1 U9275 ( .A1(n8257), .A2(n8256), .ZN(n8277) );
  NAND2_X1 U9276 ( .A1(n8464), .A2(n8631), .ZN(n8467) );
  NAND2_X1 U9277 ( .A1(n6685), .A2(n6684), .ZN(n12251) );
  INV_X1 U9278 ( .A(n12347), .ZN(n6693) );
  CLKBUF_X2 U9279 ( .A(n14265), .Z(n6688) );
  NAND2_X1 U9280 ( .A1(n9389), .A2(n12131), .ZN(n9390) );
  NAND2_X1 U9281 ( .A1(n6694), .A2(n6693), .ZN(n6692) );
  NAND2_X1 U9282 ( .A1(n6697), .A2(n6696), .ZN(n6695) );
  NAND2_X2 U9283 ( .A1(n10956), .A2(n10955), .ZN(n12514) );
  OAI21_X2 U9284 ( .B1(n9774), .B2(n12954), .A(n9777), .ZN(n10055) );
  NAND3_X1 U9285 ( .A1(n7317), .A2(n7318), .A3(n8235), .ZN(n8239) );
  NAND2_X2 U9286 ( .A1(n11072), .A2(n11087), .ZN(n11675) );
  NAND2_X1 U9287 ( .A1(n12349), .A2(n12348), .ZN(n6694) );
  NAND2_X1 U9288 ( .A1(n12217), .A2(n12216), .ZN(n6697) );
  NAND2_X1 U9289 ( .A1(n14142), .A2(n14141), .ZN(n14140) );
  NAND2_X1 U9290 ( .A1(n6860), .A2(n6858), .ZN(n14185) );
  AOI21_X1 U9291 ( .B1(n12318), .B2(n12317), .A(n12315), .ZN(n12316) );
  NAND2_X1 U9292 ( .A1(n7748), .A2(n7747), .ZN(n7543) );
  NAND2_X1 U9293 ( .A1(n7733), .A2(n7732), .ZN(n6700) );
  NAND2_X1 U9294 ( .A1(n6893), .A2(n6713), .ZN(n6715) );
  NOR2_X1 U9295 ( .A1(n13134), .A2(n6714), .ZN(n6713) );
  OAI211_X1 U9296 ( .C1(n6890), .C2(n6714), .A(n6716), .B(n6715), .ZN(n11661)
         );
  OAI21_X1 U9297 ( .B1(n6892), .B2(n13134), .A(n6890), .ZN(n13108) );
  NAND2_X1 U9298 ( .A1(n7653), .A2(n6557), .ZN(n6720) );
  NAND2_X1 U9299 ( .A1(n7576), .A2(n6720), .ZN(n7957) );
  NAND2_X1 U9300 ( .A1(n7653), .A2(n7574), .ZN(n7575) );
  NAND2_X1 U9301 ( .A1(n7580), .A2(n6721), .ZN(n7583) );
  NAND2_X1 U9302 ( .A1(n7580), .A2(n7579), .ZN(n7581) );
  INV_X1 U9303 ( .A(n7582), .ZN(n6723) );
  OAI21_X1 U9304 ( .B1(n6723), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n7583), .ZN(
        n8004) );
  NOR2_X1 U9305 ( .A1(n14709), .A2(n7497), .ZN(n7499) );
  NOR2_X1 U9306 ( .A1(n7497), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6729) );
  INV_X1 U9307 ( .A(n14709), .ZN(n6730) );
  NAND2_X1 U9308 ( .A1(n14712), .A2(n6524), .ZN(n6734) );
  AOI21_X1 U9309 ( .B1(n7523), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n6747), .ZN(
        n6738) );
  NAND2_X1 U9310 ( .A1(n14754), .A2(n6745), .ZN(n6744) );
  NAND2_X1 U9311 ( .A1(n14754), .A2(n14753), .ZN(n14752) );
  MUX2_X1 U9312 ( .A(n9171), .B(P3_REG2_REG_2__SCAN_IN), .S(n9207), .Z(n9201)
         );
  XNOR2_X2 U9313 ( .A(n7717), .B(P3_IR_REG_2__SCAN_IN), .ZN(n9207) );
  NAND2_X1 U9315 ( .A1(n13448), .A2(n6766), .ZN(n6760) );
  NAND2_X2 U9316 ( .A1(n7325), .A2(n8631), .ZN(n8834) );
  NAND2_X2 U9317 ( .A1(n13480), .A2(n7238), .ZN(n7234) );
  INV_X1 U9318 ( .A(n6769), .ZN(n6768) );
  OAI21_X1 U9319 ( .B1(n10207), .B2(n6449), .A(n10232), .ZN(n6769) );
  NAND2_X1 U9320 ( .A1(n8968), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6770) );
  NAND2_X2 U9321 ( .A1(P2_U3088), .A2(n11907), .ZN(n14088) );
  MUX2_X1 U9322 ( .A(n8840), .B(n8835), .S(n6772), .Z(n9030) );
  MUX2_X1 U9323 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6772), .Z(n9409) );
  MUX2_X1 U9324 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n6772), .Z(n10079) );
  MUX2_X1 U9325 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n6772), .Z(n10199) );
  MUX2_X1 U9326 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n6772), .Z(n10800) );
  MUX2_X1 U9327 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n6772), .Z(n11325) );
  MUX2_X1 U9328 ( .A(n14081), .B(n14681), .S(n6772), .Z(n11295) );
  NAND2_X1 U9329 ( .A1(n14456), .A2(n6776), .ZN(n6775) );
  OAI21_X1 U9330 ( .B1(n14535), .B2(n6784), .A(n6783), .ZN(n14479) );
  NAND2_X1 U9331 ( .A1(n10392), .A2(n6790), .ZN(n10526) );
  INV_X2 U9332 ( .A(n9924), .ZN(n11913) );
  NOR2_X4 U9333 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n8336) );
  INV_X2 U9334 ( .A(n11391), .ZN(n12116) );
  NOR2_X2 U9335 ( .A1(n10399), .A2(n14962), .ZN(n6800) );
  NOR2_X2 U9336 ( .A1(n14462), .A2(n14470), .ZN(n14465) );
  NOR2_X2 U9337 ( .A1(n14519), .A2(n14636), .ZN(n6802) );
  NOR2_X2 U9338 ( .A1(n14400), .A2(n14586), .ZN(n11457) );
  NOR2_X2 U9339 ( .A1(n14432), .A2(n14420), .ZN(n14419) );
  NAND2_X1 U9340 ( .A1(n14348), .A2(n6805), .ZN(n14330) );
  NAND2_X1 U9341 ( .A1(n14348), .A2(n6803), .ZN(n14337) );
  NAND2_X1 U9342 ( .A1(n14348), .A2(n12096), .ZN(n11770) );
  INV_X1 U9343 ( .A(n14330), .ZN(n14338) );
  NOR2_X2 U9344 ( .A1(n14711), .A2(n14710), .ZN(n14709) );
  XNOR2_X2 U9345 ( .A(n7503), .B(n6808), .ZN(n14713) );
  XNOR2_X1 U9346 ( .A(n9227), .B(n9226), .ZN(n14130) );
  OAI22_X2 U9347 ( .A1(n14176), .A2(n6827), .B1(n6829), .B2(n11815), .ZN(
        n14142) );
  NAND2_X1 U9348 ( .A1(n14157), .A2(n7362), .ZN(n6841) );
  OAI211_X1 U9349 ( .C1(n14157), .C2(n6839), .A(n6836), .B(n6833), .ZN(n11893)
         );
  NAND2_X1 U9350 ( .A1(n14157), .A2(n6834), .ZN(n6833) );
  OR2_X1 U9351 ( .A1(n6840), .A2(n6845), .ZN(n6837) );
  NAND2_X1 U9352 ( .A1(n6840), .A2(n6523), .ZN(n6838) );
  NAND2_X1 U9353 ( .A1(n9615), .A2(n6850), .ZN(n6849) );
  NAND2_X1 U9354 ( .A1(n11785), .A2(n6855), .ZN(n6857) );
  INV_X1 U9355 ( .A(n6857), .ZN(n14109) );
  NAND2_X1 U9356 ( .A1(n14194), .A2(n6861), .ZN(n6860) );
  INV_X2 U9357 ( .A(n11404), .ZN(n11366) );
  AND3_X2 U9358 ( .A1(n6869), .A2(n6868), .A3(n6867), .ZN(n7773) );
  NAND3_X1 U9359 ( .A1(n7417), .A2(n7894), .A3(n11095), .ZN(n6871) );
  NAND3_X1 U9360 ( .A1(n6871), .A2(n6870), .A3(n7923), .ZN(n7924) );
  NAND2_X1 U9361 ( .A1(n13183), .A2(n6883), .ZN(n6881) );
  INV_X1 U9362 ( .A(n6879), .ZN(n6886) );
  OAI22_X1 U9363 ( .A1(n7749), .A2(n8267), .B1(n9135), .B2(n9173), .ZN(n6889)
         );
  INV_X1 U9364 ( .A(n9779), .ZN(n15187) );
  NAND2_X1 U9365 ( .A1(n15173), .A2(n15187), .ZN(n12770) );
  NAND2_X1 U9366 ( .A1(n13232), .A2(n6897), .ZN(n6895) );
  NAND2_X1 U9367 ( .A1(n6896), .A2(n6895), .ZN(n13199) );
  NAND2_X1 U9368 ( .A1(n10578), .A2(n7798), .ZN(n6912) );
  AND2_X1 U9369 ( .A1(n6912), .A2(n7796), .ZN(n10814) );
  NAND2_X1 U9370 ( .A1(n11158), .A2(n11157), .ZN(n6914) );
  NAND2_X1 U9371 ( .A1(n11158), .A2(n6920), .ZN(n6915) );
  NAND2_X1 U9372 ( .A1(n8834), .A2(n6938), .ZN(n6935) );
  NAND2_X2 U9373 ( .A1(n8500), .A2(n8606), .ZN(n8931) );
  NOR2_X2 U9374 ( .A1(n13879), .A2(n14050), .ZN(n13842) );
  NOR2_X2 U9375 ( .A1(n10252), .A2(n6651), .ZN(n10363) );
  NAND2_X1 U9376 ( .A1(n11627), .A2(n6952), .ZN(n13775) );
  INV_X1 U9377 ( .A(n14076), .ZN(n6960) );
  AND2_X4 U9378 ( .A1(n14073), .A2(n6960), .ZN(n12390) );
  INV_X1 U9379 ( .A(n8680), .ZN(n12447) );
  NAND2_X1 U9380 ( .A1(n9732), .A2(n8680), .ZN(n8842) );
  OAI211_X2 U9381 ( .C1(n8931), .C2(n8672), .A(n8671), .B(n8670), .ZN(n13926)
         );
  INV_X1 U9382 ( .A(n8585), .ZN(n8587) );
  OAI21_X1 U9383 ( .B1(n6964), .B2(n14068), .A(P2_IR_REG_29__SCAN_IN), .ZN(
        n6963) );
  NAND2_X1 U9384 ( .A1(n13792), .A2(n6968), .ZN(n6966) );
  OAI21_X1 U9385 ( .B1(n13840), .B2(n6982), .A(n6980), .ZN(n13802) );
  INV_X1 U9386 ( .A(n13840), .ZN(n6986) );
  NAND2_X1 U9387 ( .A1(n6991), .A2(n12466), .ZN(n6989) );
  NAND2_X1 U9388 ( .A1(n11634), .A2(n6451), .ZN(n6998) );
  NAND2_X1 U9389 ( .A1(n10921), .A2(n7003), .ZN(n7002) );
  NAND2_X1 U9390 ( .A1(n7009), .A2(n7008), .ZN(P3_U3296) );
  NAND2_X1 U9391 ( .A1(n7010), .A2(n12963), .ZN(n7009) );
  NAND2_X1 U9392 ( .A1(n7011), .A2(n12958), .ZN(n7010) );
  NAND2_X1 U9393 ( .A1(n7012), .A2(n12761), .ZN(n7011) );
  XNOR2_X1 U9394 ( .A(n12760), .B(n13072), .ZN(n7012) );
  NAND2_X1 U9395 ( .A1(n7016), .A2(n7013), .ZN(n13147) );
  NAND3_X1 U9396 ( .A1(n13189), .A2(n7017), .A3(n6471), .ZN(n7016) );
  NAND2_X1 U9397 ( .A1(n10597), .A2(n7024), .ZN(n7023) );
  AOI21_X1 U9398 ( .B1(n7024), .B2(n7026), .A(n7022), .ZN(n7021) );
  INV_X1 U9399 ( .A(n12812), .ZN(n7022) );
  NAND2_X1 U9400 ( .A1(n14757), .A2(n7030), .ZN(n7028) );
  INV_X1 U9401 ( .A(n7037), .ZN(n12759) );
  AOI21_X1 U9402 ( .B1(n11655), .B2(n6462), .A(n6429), .ZN(n7040) );
  AOI21_X1 U9403 ( .B1(n11655), .B2(n12947), .A(n12902), .ZN(n13086) );
  NAND2_X1 U9404 ( .A1(n13146), .A2(n6528), .ZN(n7056) );
  CLKBUF_X1 U9405 ( .A(n7056), .Z(n7054) );
  NAND2_X1 U9406 ( .A1(n13146), .A2(n12763), .ZN(n13139) );
  NAND2_X1 U9407 ( .A1(n7603), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7602) );
  AND2_X1 U9408 ( .A1(n7682), .A2(n7058), .ZN(n7057) );
  NOR2_X2 U9409 ( .A1(n8163), .A2(n8162), .ZN(n8181) );
  NOR2_X2 U9410 ( .A1(n7079), .A2(n7080), .ZN(n9422) );
  OAI22_X1 U9411 ( .A1(n13854), .A2(n11535), .B1(n13541), .B2(n14050), .ZN(
        n13840) );
  NAND2_X1 U9412 ( .A1(n10240), .A2(n10239), .ZN(n10369) );
  NAND2_X1 U9413 ( .A1(n13606), .A2(n13605), .ZN(n13607) );
  NAND2_X1 U9414 ( .A1(n8876), .A2(n8875), .ZN(n8874) );
  AND2_X2 U9415 ( .A1(n9395), .A2(n11936), .ZN(n9519) );
  NAND2_X1 U9416 ( .A1(n7078), .A2(n8181), .ZN(n8325) );
  NOR2_X2 U9417 ( .A1(n9518), .A2(n14135), .ZN(n9509) );
  NOR2_X2 U9418 ( .A1(n10009), .A2(n14096), .ZN(n10271) );
  NOR2_X2 U9419 ( .A1(n10319), .A2(n15097), .ZN(n10318) );
  NOR2_X2 U9420 ( .A1(n13580), .A2(n13777), .ZN(n13934) );
  NOR2_X2 U9421 ( .A1(n8878), .A2(n13908), .ZN(n10292) );
  NOR2_X2 U9422 ( .A1(n13944), .A2(n13601), .ZN(n13586) );
  AOI21_X1 U9423 ( .B1(n7063), .B2(n8990), .A(n7062), .ZN(n7064) );
  NOR2_X1 U9424 ( .A1(n11404), .A2(n7065), .ZN(n7062) );
  INV_X1 U9425 ( .A(n9924), .ZN(n7063) );
  NAND2_X2 U9426 ( .A1(n11404), .A2(n8968), .ZN(n9924) );
  AND2_X2 U9427 ( .A1(n7064), .A2(n8992), .ZN(n14933) );
  INV_X1 U9428 ( .A(n8991), .ZN(n7065) );
  OAI21_X1 U9429 ( .B1(n14360), .B2(n7072), .A(n7070), .ZN(n7073) );
  INV_X1 U9430 ( .A(n8336), .ZN(n7079) );
  OAI21_X1 U9431 ( .B1(n7084), .B2(n9685), .A(n7082), .ZN(n9942) );
  AOI21_X1 U9432 ( .B1(n7086), .B2(n7083), .A(n7085), .ZN(n7082) );
  INV_X1 U9433 ( .A(n7086), .ZN(n7084) );
  NAND2_X1 U9434 ( .A1(n11955), .A2(n7097), .ZN(n11960) );
  INV_X1 U9435 ( .A(n11958), .ZN(n7097) );
  NAND2_X1 U9436 ( .A1(n7321), .A2(n6473), .ZN(n7098) );
  NAND2_X1 U9437 ( .A1(n12101), .A2(n12102), .ZN(n7113) );
  NAND2_X1 U9438 ( .A1(n7115), .A2(n7116), .ZN(n7114) );
  NAND2_X1 U9439 ( .A1(n12100), .A2(n12099), .ZN(n7115) );
  NAND2_X1 U9440 ( .A1(n12095), .A2(n12094), .ZN(n12100) );
  INV_X1 U9441 ( .A(n11996), .ZN(n7119) );
  NAND3_X1 U9442 ( .A1(n12084), .A2(n12083), .A3(n6534), .ZN(n7121) );
  INV_X1 U9443 ( .A(n12085), .ZN(n7122) );
  NAND2_X1 U9444 ( .A1(n11976), .A2(n7123), .ZN(n7127) );
  NAND2_X1 U9445 ( .A1(n8167), .A2(n7135), .ZN(n8320) );
  NAND2_X1 U9446 ( .A1(n7142), .A2(n7144), .ZN(n12032) );
  NAND3_X1 U9447 ( .A1(n12013), .A2(n12012), .A3(n7143), .ZN(n7142) );
  AOI21_X1 U9448 ( .B1(n12019), .B2(n12014), .A(n6510), .ZN(n7144) );
  NAND3_X1 U9449 ( .A1(n7168), .A2(n7167), .A3(n7166), .ZN(n7165) );
  OAI21_X2 U9450 ( .B1(n7994), .B2(n7172), .A(n7169), .ZN(n8015) );
  INV_X1 U9451 ( .A(n7170), .ZN(n7169) );
  NAND2_X1 U9452 ( .A1(n11649), .A2(n7175), .ZN(n7173) );
  OAI21_X1 U9453 ( .B1(n13772), .B2(n7189), .A(n7184), .ZN(n13591) );
  NAND2_X1 U9454 ( .A1(n9765), .A2(n6430), .ZN(n7194) );
  NAND2_X1 U9455 ( .A1(n13835), .A2(n7201), .ZN(n7200) );
  NAND2_X1 U9456 ( .A1(n10312), .A2(n7208), .ZN(n7207) );
  NAND2_X1 U9457 ( .A1(n9593), .A2(n7212), .ZN(n8493) );
  MUX2_X1 U9458 ( .A(n13950), .B(n7215), .S(n15112), .Z(n13951) );
  MUX2_X1 U9459 ( .A(n14030), .B(n7215), .S(n15106), .Z(n14031) );
  NAND2_X1 U9460 ( .A1(n13873), .A2(n13877), .ZN(n7219) );
  NAND2_X1 U9462 ( .A1(n7234), .A2(n7235), .ZN(n13458) );
  OAI21_X1 U9463 ( .B1(n9697), .B2(n9696), .A(n9702), .ZN(n9720) );
  INV_X1 U9464 ( .A(n7249), .ZN(n14371) );
  INV_X1 U9465 ( .A(n9395), .ZN(n14920) );
  XNOR2_X2 U9466 ( .A(n14265), .B(n9395), .ZN(n12131) );
  AND3_X2 U9467 ( .A1(n8971), .A2(n8970), .A3(n6470), .ZN(n9395) );
  NAND2_X1 U9468 ( .A1(n11177), .A2(n6530), .ZN(n11183) );
  NAND2_X1 U9469 ( .A1(n14458), .A2(n7251), .ZN(n7250) );
  NAND2_X1 U9470 ( .A1(n7250), .A2(n7253), .ZN(n14411) );
  NAND2_X1 U9471 ( .A1(n7264), .A2(n7263), .ZN(n11365) );
  AND2_X1 U9472 ( .A1(n11445), .A2(n7265), .ZN(n7263) );
  INV_X1 U9473 ( .A(n10057), .ZN(n7277) );
  NAND2_X1 U9474 ( .A1(n7295), .A2(n7293), .ZN(n10671) );
  OAI21_X2 U9475 ( .B1(n12672), .B2(n7300), .A(n7298), .ZN(n12550) );
  OAI21_X2 U9476 ( .B1(n12514), .B2(n7305), .A(n7303), .ZN(n12683) );
  NAND2_X1 U9477 ( .A1(n7654), .A2(n6432), .ZN(n8029) );
  INV_X1 U9478 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7314) );
  INV_X1 U9479 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7316) );
  NAND3_X1 U9480 ( .A1(n8231), .A2(n8233), .A3(n8230), .ZN(n7317) );
  INV_X1 U9481 ( .A(n8239), .ZN(n8253) );
  NAND2_X1 U9482 ( .A1(n12107), .A2(n12106), .ZN(n7322) );
  NAND2_X1 U9483 ( .A1(n12108), .A2(n12109), .ZN(n7323) );
  NAND2_X1 U9484 ( .A1(n10078), .A2(n7329), .ZN(n7328) );
  INV_X1 U9485 ( .A(n11331), .ZN(n7343) );
  NAND2_X1 U9486 ( .A1(n10798), .A2(n10745), .ZN(n11402) );
  INV_X1 U9487 ( .A(n10747), .ZN(n7352) );
  NAND2_X4 U9488 ( .A1(n8695), .A2(n7356), .ZN(n11919) );
  NAND3_X1 U9489 ( .A1(n8326), .A2(n7377), .A3(n8327), .ZN(n7376) );
  NAND2_X1 U9490 ( .A1(n9216), .A2(n7378), .ZN(n14132) );
  NAND3_X2 U9491 ( .A1(n10750), .A2(n12488), .A3(n12489), .ZN(n12432) );
  NAND2_X1 U9492 ( .A1(n13561), .A2(n12223), .ZN(n12191) );
  NAND2_X1 U9493 ( .A1(n8587), .A2(n7384), .ZN(n8591) );
  INV_X1 U9494 ( .A(n12304), .ZN(n7386) );
  INV_X1 U9495 ( .A(n12305), .ZN(n7387) );
  NAND3_X1 U9496 ( .A1(n12239), .A2(n6536), .A3(n12238), .ZN(n7388) );
  INV_X1 U9497 ( .A(n12333), .ZN(n7392) );
  NAND2_X1 U9498 ( .A1(n7393), .A2(n7394), .ZN(n12277) );
  NAND2_X1 U9499 ( .A1(n10688), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8677) );
  MUX2_X2 U9500 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n8127), .S(n15232), .Z(n8128) );
  MUX2_X2 U9501 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n8127), .S(n15240), .Z(n8114) );
  MUX2_X1 U9502 ( .A(n14920), .B(n6688), .S(n11933), .Z(n11942) );
  XNOR2_X1 U9503 ( .A(n11614), .B(n7007), .ZN(n11626) );
  OAI22_X1 U9504 ( .A1(n10851), .A2(n10850), .B1(n10849), .B2(n14256), .ZN(
        n14725) );
  OAI21_X1 U9506 ( .B1(n7614), .B2(n7613), .A(P3_IR_REG_29__SCAN_IN), .ZN(
        n7616) );
  NAND2_X1 U9507 ( .A1(n7614), .A2(n7610), .ZN(n7612) );
  NAND2_X1 U9508 ( .A1(n8493), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8494) );
  AND2_X4 U9509 ( .A1(n12506), .A2(n13397), .ZN(n7852) );
  NAND2_X1 U9510 ( .A1(n8074), .A2(n8073), .ZN(n8084) );
  NAND2_X1 U9511 ( .A1(n12770), .A2(n15190), .ZN(n9782) );
  NAND2_X1 U9512 ( .A1(n11288), .A2(n6918), .ZN(n11331) );
  AND3_X2 U9513 ( .A1(n7709), .A2(n7708), .A3(n7707), .ZN(n12771) );
  INV_X1 U9514 ( .A(n8242), .ZN(n8244) );
  AND2_X1 U9515 ( .A1(n9248), .A2(n8348), .ZN(n8805) );
  NAND2_X4 U9516 ( .A1(n8696), .A2(n8693), .ZN(n9229) );
  NAND2_X1 U9517 ( .A1(n8236), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8205) );
  AND3_X1 U9518 ( .A1(n6667), .A2(n12179), .A3(n12443), .ZN(n15098) );
  INV_X1 U9519 ( .A(n14073), .ZN(n8593) );
  AND2_X1 U9520 ( .A1(n15101), .A2(n12181), .ZN(n12186) );
  AND2_X1 U9521 ( .A1(n6597), .A2(n15101), .ZN(n15093) );
  OR2_X1 U9522 ( .A1(n15101), .A2(n12441), .ZN(n9099) );
  NOR2_X1 U9523 ( .A1(n7850), .A2(n7849), .ZN(n7402) );
  AND2_X1 U9524 ( .A1(n12756), .A2(n13081), .ZN(n7404) );
  AND2_X1 U9525 ( .A1(n12753), .A2(n12912), .ZN(n7405) );
  NAND2_X1 U9526 ( .A1(n9128), .A2(n13825), .ZN(n13868) );
  AND2_X1 U9527 ( .A1(n9610), .A2(n9611), .ZN(n7406) );
  AND2_X1 U9528 ( .A1(n11667), .A2(n7422), .ZN(n7407) );
  OR2_X1 U9529 ( .A1(n13101), .A2(n13384), .ZN(n7408) );
  OR2_X1 U9530 ( .A1(n13101), .A2(n13334), .ZN(n7409) );
  AND2_X1 U9531 ( .A1(n14489), .A2(n14494), .ZN(n7410) );
  OR2_X1 U9532 ( .A1(n11723), .A2(n11722), .ZN(n7411) );
  OR2_X1 U9533 ( .A1(n13289), .A2(n12644), .ZN(n7412) );
  AND2_X1 U9534 ( .A1(n6688), .A2(n9395), .ZN(n7414) );
  AND2_X1 U9535 ( .A1(n9783), .A2(n9782), .ZN(n7416) );
  AND2_X1 U9536 ( .A1(n7908), .A2(n7418), .ZN(n7417) );
  OR2_X1 U9537 ( .A1(n13385), .A2(n13247), .ZN(n7418) );
  AND2_X1 U9538 ( .A1(n13610), .A2(n13609), .ZN(n7419) );
  OR2_X1 U9539 ( .A1(n14265), .A2(n14920), .ZN(n7420) );
  INV_X1 U9540 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10426) );
  OR2_X1 U9541 ( .A1(n12755), .A2(n13080), .ZN(n7422) );
  AND2_X1 U9542 ( .A1(n12379), .A2(n12368), .ZN(n7423) );
  INV_X2 U9543 ( .A(n15241), .ZN(n15240) );
  XNOR2_X1 U9544 ( .A(n14334), .B(n12159), .ZN(n7424) );
  INV_X1 U9545 ( .A(n12139), .ZN(n10545) );
  OR2_X1 U9546 ( .A1(n12124), .A2(n11936), .ZN(n11939) );
  OR2_X1 U9547 ( .A1(n11971), .A2(n11970), .ZN(n11976) );
  INV_X1 U9548 ( .A(n12246), .ZN(n12247) );
  INV_X1 U9549 ( .A(n12071), .ZN(n12072) );
  OR2_X1 U9550 ( .A1(n12373), .A2(n12372), .ZN(n12368) );
  MUX2_X1 U9551 ( .A(n12097), .B(n12096), .S(n12119), .Z(n12098) );
  INV_X1 U9552 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7595) );
  INV_X1 U9553 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8160) );
  OR2_X1 U9554 ( .A1(n12736), .A2(n13263), .ZN(n7923) );
  INV_X1 U9555 ( .A(n12430), .ZN(n12417) );
  INV_X1 U9556 ( .A(n13855), .ZN(n11535) );
  INV_X1 U9557 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8143) );
  INV_X1 U9558 ( .A(n12138), .ZN(n10277) );
  NOR2_X1 U9559 ( .A1(n12757), .A2(n7404), .ZN(n12758) );
  INV_X1 U9560 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n12651) );
  INV_X1 U9561 ( .A(n11075), .ZN(n11073) );
  INV_X1 U9562 ( .A(n11555), .ZN(n11478) );
  INV_X1 U9563 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10840) );
  INV_X1 U9564 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n14112) );
  INV_X1 U9565 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9417) );
  INV_X1 U9566 ( .A(n10959), .ZN(n10955) );
  OR2_X1 U9567 ( .A1(n7975), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n7977) );
  NAND2_X1 U9568 ( .A1(n7924), .A2(n7413), .ZN(n13232) );
  INV_X1 U9569 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n7799) );
  INV_X1 U9570 ( .A(n14772), .ZN(n8056) );
  AND2_X1 U9571 ( .A1(n7557), .A2(n7556), .ZN(n7864) );
  INV_X1 U9572 ( .A(n13506), .ZN(n11680) );
  INV_X1 U9573 ( .A(n12181), .ZN(n12444) );
  OR2_X1 U9574 ( .A1(n11582), .A2(n11493), .ZN(n11592) );
  OR2_X1 U9575 ( .A1(n11542), .A2(n11477), .ZN(n11555) );
  NAND2_X1 U9576 ( .A1(n11073), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n11233) );
  INV_X1 U9577 ( .A(n13604), .ZN(n13605) );
  NAND2_X1 U9578 ( .A1(n11478), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n11569) );
  OR2_X1 U9579 ( .A1(n9859), .A2(n9858), .ZN(n10214) );
  NAND2_X1 U9580 ( .A1(n12448), .A2(n8866), .ZN(n10300) );
  INV_X1 U9581 ( .A(n13574), .ZN(n8602) );
  XNOR2_X1 U9582 ( .A(n6667), .B(n12181), .ZN(n8605) );
  AOI21_X1 U9583 ( .B1(n8572), .B2(n8571), .A(n8570), .ZN(n9089) );
  NAND2_X1 U9584 ( .A1(n8153), .A2(n8152), .ZN(n8155) );
  OR2_X1 U9585 ( .A1(n9546), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n9042) );
  INV_X1 U9586 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8137) );
  OR2_X1 U9587 ( .A1(n11025), .A2(n11024), .ZN(n11026) );
  INV_X1 U9588 ( .A(n14168), .ZN(n11799) );
  NAND2_X1 U9589 ( .A1(n11407), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11406) );
  INV_X1 U9590 ( .A(n12170), .ZN(n12171) );
  NAND2_X1 U9591 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n11345), .ZN(n11344) );
  NAND2_X1 U9592 ( .A1(n11303), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11434) );
  INV_X1 U9593 ( .A(n12133), .ZN(n10014) );
  INV_X1 U9594 ( .A(n14243), .ZN(n11887) );
  OR2_X1 U9595 ( .A1(n11164), .A2(P1_B_REG_SCAN_IN), .ZN(n8344) );
  INV_X1 U9596 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8166) );
  OR2_X1 U9597 ( .A1(n8827), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8828) );
  INV_X1 U9598 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7445) );
  INV_X1 U9599 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n13709) );
  OR2_X1 U9600 ( .A1(n7673), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7962) );
  INV_X1 U9601 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9379) );
  OR2_X1 U9602 ( .A1(n7996), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8008) );
  NAND2_X1 U9603 ( .A1(n7625), .A2(n7624), .ZN(n7975) );
  OR2_X1 U9604 ( .A1(n9787), .A2(n9674), .ZN(n12734) );
  AND4_X1 U9605 ( .A1(n10039), .A2(n10038), .A3(n10037), .A4(n10036), .ZN(
        n13089) );
  INV_X1 U9606 ( .A(n10789), .ZN(n10767) );
  AND2_X1 U9607 ( .A1(n9144), .A2(n9142), .ZN(n9139) );
  INV_X1 U9608 ( .A(n12926), .ZN(n13124) );
  INV_X1 U9609 ( .A(n13200), .ZN(n13174) );
  AND2_X2 U9610 ( .A1(n9830), .A2(n12773), .ZN(n12917) );
  INV_X1 U9611 ( .A(n14759), .ZN(n13247) );
  NAND2_X1 U9612 ( .A1(n9661), .A2(n13387), .ZN(n9672) );
  INV_X1 U9613 ( .A(n9776), .ZN(n13072) );
  AND2_X1 U9614 ( .A1(n13386), .A2(n13388), .ZN(n8116) );
  INV_X1 U9615 ( .A(n12968), .ZN(n12700) );
  AND2_X1 U9616 ( .A1(n7566), .A2(n7565), .ZN(n7909) );
  AND2_X1 U9617 ( .A1(n7551), .A2(n7550), .ZN(n7811) );
  AND2_X1 U9618 ( .A1(n7542), .A2(n7541), .ZN(n7747) );
  INV_X1 U9619 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n11084) );
  OR2_X1 U9620 ( .A1(n10220), .A2(n10426), .ZN(n10418) );
  OR2_X1 U9621 ( .A1(n9089), .A2(n9086), .ZN(n9101) );
  AND2_X1 U9622 ( .A1(n11592), .A2(n11494), .ZN(n13778) );
  OR2_X1 U9623 ( .A1(n10418), .A2(n11706), .ZN(n10654) );
  INV_X1 U9624 ( .A(n8522), .ZN(n8521) );
  NAND2_X1 U9625 ( .A1(n13582), .A2(n13532), .ZN(n11623) );
  INV_X1 U9626 ( .A(n13891), .ZN(n13875) );
  AND2_X1 U9627 ( .A1(n14089), .A2(n8568), .ZN(n8569) );
  NAND2_X1 U9628 ( .A1(n8155), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8142) );
  OR2_X1 U9629 ( .A1(n11801), .A2(n11800), .ZN(n11802) );
  OR2_X1 U9630 ( .A1(n8807), .A2(n14540), .ZN(n8808) );
  INV_X1 U9631 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10116) );
  OR2_X1 U9632 ( .A1(n11927), .A2(n8764), .ZN(n9249) );
  OR2_X1 U9633 ( .A1(n14233), .A2(n14637), .ZN(n14871) );
  OR2_X1 U9634 ( .A1(n9247), .A2(n9265), .ZN(n14233) );
  AND2_X1 U9635 ( .A1(n14296), .A2(n11051), .ZN(n14308) );
  INV_X1 U9636 ( .A(n14566), .ZN(n12096) );
  INV_X1 U9637 ( .A(n12147), .ZN(n10972) );
  INV_X1 U9638 ( .A(n12136), .ZN(n9944) );
  INV_X1 U9639 ( .A(n6699), .ZN(n11930) );
  OR2_X1 U9640 ( .A1(n9268), .A2(n11367), .ZN(n14497) );
  XNOR2_X1 U9641 ( .A(n10079), .B(n10080), .ZN(n10077) );
  AOI22_X1 U9642 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n7439), .B1(n7495), .B2(
        n7438), .ZN(n7441) );
  OAI21_X1 U9643 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n13709), .A(n7457), .ZN(
        n7469) );
  NAND2_X1 U9644 ( .A1(n9670), .A2(n9669), .ZN(n12729) );
  XNOR2_X1 U9645 ( .A(n8031), .B(n8030), .ZN(n12962) );
  AND4_X1 U9646 ( .A1(n8043), .A2(n8042), .A3(n8041), .A4(n8040), .ZN(n12569)
         );
  AND4_X1 U9647 ( .A1(n7991), .A2(n7990), .A3(n7989), .A4(n7988), .ZN(n13164)
         );
  INV_X1 U9648 ( .A(n15140), .ZN(n13023) );
  AND2_X1 U9649 ( .A1(n9139), .A2(n9138), .ZN(n15154) );
  AND3_X1 U9650 ( .A1(n9137), .A2(n12917), .A3(n9135), .ZN(n15192) );
  INV_X1 U9651 ( .A(n13207), .ZN(n13270) );
  INV_X1 U9652 ( .A(n15169), .ZN(n15201) );
  OR3_X1 U9653 ( .A1(n8116), .A2(n8107), .A3(n8106), .ZN(n9792) );
  INV_X1 U9654 ( .A(n15226), .ZN(n13311) );
  AND2_X1 U9655 ( .A1(n15177), .A2(n15228), .ZN(n14790) );
  INV_X1 U9656 ( .A(n14790), .ZN(n14798) );
  INV_X1 U9657 ( .A(n15228), .ZN(n15223) );
  INV_X1 U9658 ( .A(n12962), .ZN(n9830) );
  NAND2_X1 U9659 ( .A1(n7883), .A2(n7882), .ZN(n7885) );
  INV_X1 U9660 ( .A(n13503), .ZN(n13521) );
  OR2_X1 U9661 ( .A1(n13602), .A2(n11606), .ZN(n11487) );
  INV_X1 U9662 ( .A(n12390), .ZN(n11609) );
  INV_X1 U9663 ( .A(n6638), .ZN(n11606) );
  NAND2_X1 U9664 ( .A1(n8521), .A2(n8503), .ZN(n15046) );
  INV_X1 U9665 ( .A(n15046), .ZN(n15003) );
  NAND2_X1 U9666 ( .A1(n8604), .A2(n8603), .ZN(n13891) );
  INV_X1 U9667 ( .A(n13871), .ZN(n15072) );
  INV_X1 U9668 ( .A(n14064), .ZN(n14051) );
  NOR2_X1 U9669 ( .A1(n14084), .A2(n8569), .ZN(n15076) );
  NOR2_X1 U9670 ( .A1(n9043), .A2(n9407), .ZN(n15051) );
  INV_X1 U9671 ( .A(n14871), .ZN(n14217) );
  INV_X1 U9672 ( .A(n14883), .ZN(n14236) );
  AND4_X1 U9673 ( .A1(n11412), .A2(n11411), .A3(n11410), .A4(n11409), .ZN(
        n14150) );
  INV_X1 U9674 ( .A(n14906), .ZN(n14318) );
  INV_X1 U9675 ( .A(n14924), .ZN(n14736) );
  NAND2_X1 U9676 ( .A1(n11761), .A2(n11760), .ZN(n11762) );
  NOR2_X1 U9677 ( .A1(n14743), .A2(n14724), .ZN(n14480) );
  INV_X1 U9678 ( .A(n14497), .ZN(n14729) );
  INV_X1 U9679 ( .A(n14506), .ZN(n14733) );
  NAND2_X1 U9680 ( .A1(n11466), .A2(n14541), .ZN(n14544) );
  INV_X1 U9681 ( .A(n9460), .ZN(n8781) );
  INV_X1 U9682 ( .A(n14832), .ZN(n14724) );
  OR2_X1 U9683 ( .A1(n11916), .A2(n11930), .ZN(n14966) );
  AOI21_X1 U9684 ( .B1(n8780), .B2(n8779), .A(n8778), .ZN(n9459) );
  XNOR2_X1 U9685 ( .A(n8186), .B(n8185), .ZN(n8330) );
  AND2_X1 U9686 ( .A1(n9426), .A2(n9534), .ZN(n14902) );
  AND2_X1 U9687 ( .A1(n8470), .A2(n8370), .ZN(n10380) );
  INV_X1 U9688 ( .A(n13387), .ZN(n8898) );
  NAND2_X1 U9689 ( .A1(n9673), .A2(n9800), .ZN(n12720) );
  NAND4_X1 U9690 ( .A1(n8024), .A2(n8023), .A3(n8022), .A4(n8021), .ZN(n13125)
         );
  INV_X1 U9691 ( .A(n13235), .ZN(n13263) );
  INV_X1 U9692 ( .A(n13071), .ZN(n15150) );
  INV_X1 U9693 ( .A(n15113), .ZN(n15157) );
  NAND2_X1 U9694 ( .A1(n9800), .A2(n15182), .ZN(n15169) );
  NAND2_X1 U9695 ( .A1(n15204), .A2(n14779), .ZN(n13207) );
  OR2_X1 U9696 ( .A1(n9792), .A2(n8113), .ZN(n15241) );
  AND2_X1 U9697 ( .A1(n14787), .A2(n14786), .ZN(n14800) );
  INV_X2 U9698 ( .A(n15234), .ZN(n15232) );
  CLKBUF_X1 U9699 ( .A(n8901), .Z(n8927) );
  INV_X1 U9700 ( .A(SI_17_), .ZN(n10080) );
  INV_X1 U9701 ( .A(SI_12_), .ZN(n9029) );
  INV_X1 U9702 ( .A(n13510), .ZN(n13525) );
  NAND2_X1 U9703 ( .A1(n9597), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13495) );
  NAND2_X1 U9704 ( .A1(n11487), .A2(n11486), .ZN(n13534) );
  INV_X1 U9705 ( .A(n14987), .ZN(n15061) );
  INV_X1 U9706 ( .A(n13927), .ZN(n15069) );
  OR2_X1 U9707 ( .A1(n15075), .A2(n9808), .ZN(n13871) );
  AND2_X2 U9708 ( .A1(n8798), .A2(n9125), .ZN(n15112) );
  INV_X1 U9709 ( .A(n13846), .ZN(n14047) );
  INV_X1 U9710 ( .A(n12300), .ZN(n10919) );
  INV_X1 U9711 ( .A(n15106), .ZN(n15104) );
  NAND2_X1 U9712 ( .A1(n15106), .A2(n15098), .ZN(n14064) );
  NOR2_X1 U9713 ( .A1(n15082), .A2(n15076), .ZN(n15080) );
  INV_X1 U9714 ( .A(n15080), .ZN(n15081) );
  INV_X1 U9715 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n13726) );
  INV_X1 U9716 ( .A(n14734), .ZN(n14745) );
  OR3_X1 U9717 ( .A1(n9247), .A2(n8810), .A3(n8809), .ZN(n14875) );
  OR2_X1 U9718 ( .A1(n14894), .A2(n9002), .ZN(n14320) );
  OR2_X1 U9719 ( .A1(n14894), .A2(n8389), .ZN(n14906) );
  INV_X1 U9720 ( .A(n14891), .ZN(n14911) );
  INV_X1 U9721 ( .A(n14739), .ZN(n14486) );
  INV_X2 U9722 ( .A(n14544), .ZN(n14743) );
  INV_X1 U9723 ( .A(n14740), .ZN(n14508) );
  AND2_X2 U9724 ( .A1(n8781), .A2(n9459), .ZN(n14986) );
  NOR2_X2 U9725 ( .A1(n9460), .A2(n9459), .ZN(n14953) );
  AND2_X1 U9726 ( .A1(n8330), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8348) );
  INV_X1 U9727 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14681) );
  INV_X1 U9728 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9588) );
  INV_X1 U9729 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8835) );
  NOR2_X2 U9730 ( .A1(n9661), .A2(n8898), .ZN(P3_U3897) );
  NAND2_X1 U9731 ( .A1(n8115), .A2(n7409), .ZN(P3_U3486) );
  NAND2_X1 U9732 ( .A1(n8129), .A2(n7408), .ZN(P3_U3454) );
  INV_X1 U9733 ( .A(n13562), .ZN(P2_U3947) );
  INV_X1 U9734 ( .A(n14266), .ZN(P1_U4016) );
  XNOR2_X1 U9735 ( .A(n7532), .B(n7531), .ZN(SUB_1596_U4) );
  XNOR2_X1 U9736 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n7525) );
  INV_X1 U9737 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7462) );
  XNOR2_X1 U9738 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7464) );
  INV_X1 U9739 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7459) );
  AND2_X1 U9740 ( .A1(n7459), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n7460) );
  INV_X1 U9741 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n13653) );
  INV_X1 U9742 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14912) );
  NAND2_X1 U9743 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14912), .ZN(n7458) );
  NOR2_X1 U9744 ( .A1(P3_ADDR_REG_14__SCAN_IN), .A2(n13709), .ZN(n7427) );
  AOI21_X1 U9745 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n13709), .A(n7427), .ZN(
        n7515) );
  INV_X1 U9746 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7456) );
  INV_X1 U9747 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n7454) );
  XNOR2_X1 U9748 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7470) );
  INV_X1 U9749 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n7452) );
  AND2_X1 U9750 ( .A1(n7452), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n7451) );
  INV_X1 U9751 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7447) );
  XNOR2_X1 U9752 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(n7447), .ZN(n7475) );
  XOR2_X1 U9753 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n7445), .Z(n7501) );
  INV_X1 U9754 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n7439) );
  NAND2_X1 U9755 ( .A1(n7481), .A2(n7480), .ZN(n7428) );
  NAND2_X1 U9756 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n7429), .ZN(n7431) );
  NAND2_X1 U9757 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n7432), .ZN(n7433) );
  NAND2_X1 U9758 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n7434), .ZN(n7437) );
  INV_X1 U9759 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7435) );
  NAND2_X1 U9760 ( .A1(n7489), .A2(n7435), .ZN(n7436) );
  NAND2_X1 U9761 ( .A1(n7437), .A2(n7436), .ZN(n7495) );
  INV_X1 U9762 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15133) );
  NAND2_X1 U9763 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n15133), .ZN(n7438) );
  INV_X1 U9764 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n7440) );
  NAND2_X1 U9765 ( .A1(n7441), .A2(n7440), .ZN(n7443) );
  XNOR2_X1 U9766 ( .A(n7441), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n7498) );
  NAND2_X1 U9767 ( .A1(n7498), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n7442) );
  NAND2_X1 U9768 ( .A1(n7443), .A2(n7442), .ZN(n7502) );
  NAND2_X1 U9769 ( .A1(n7501), .A2(n7502), .ZN(n7444) );
  NAND2_X1 U9770 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n7448), .ZN(n7450) );
  XNOR2_X1 U9771 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n7448), .ZN(n7509) );
  NAND2_X1 U9772 ( .A1(n7470), .A2(n7471), .ZN(n7453) );
  OR2_X1 U9773 ( .A1(n7456), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n7455) );
  AOI22_X1 U9774 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n7456), .B1(n7512), .B2(
        n7455), .ZN(n7514) );
  NAND2_X1 U9775 ( .A1(n7515), .A2(n7514), .ZN(n7457) );
  AOI22_X1 U9776 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n13653), .B1(n7458), .B2(
        n7469), .ZN(n7466) );
  OAI22_X1 U9777 ( .A1(n7460), .A2(n7466), .B1(P3_ADDR_REG_16__SCAN_IN), .B2(
        n7459), .ZN(n7463) );
  NAND2_X1 U9778 ( .A1(n7464), .A2(n7463), .ZN(n7461) );
  OAI21_X1 U9779 ( .B1(P3_ADDR_REG_17__SCAN_IN), .B2(n7462), .A(n7461), .ZN(
        n7524) );
  XNOR2_X1 U9780 ( .A(n7464), .B(n7463), .ZN(n7521) );
  XOR2_X1 U9781 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .Z(n7465) );
  XNOR2_X1 U9782 ( .A(n7466), .B(n7465), .ZN(n14867) );
  NAND2_X1 U9783 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n13653), .ZN(n7467) );
  OAI21_X1 U9784 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n13653), .A(n7467), .ZN(
        n7468) );
  XNOR2_X1 U9785 ( .A(n7469), .B(n7468), .ZN(n7518) );
  XOR2_X1 U9786 ( .A(n7471), .B(n7470), .Z(n14849) );
  XNOR2_X1 U9787 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7473) );
  XNOR2_X1 U9788 ( .A(n7473), .B(n7472), .ZN(n14845) );
  XOR2_X1 U9789 ( .A(n7475), .B(n7474), .Z(n7506) );
  INV_X1 U9790 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n15015) );
  NOR2_X1 U9791 ( .A1(n7487), .A2(n15015), .ZN(n7488) );
  XNOR2_X1 U9792 ( .A(n7477), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n15255) );
  XOR2_X1 U9793 ( .A(n7479), .B(n7478), .Z(n14707) );
  INV_X1 U9794 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n8650) );
  NOR2_X1 U9795 ( .A1(n7484), .A2(n8650), .ZN(n7485) );
  OAI21_X1 U9796 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n7483), .A(n7482), .ZN(
        n15249) );
  NAND2_X1 U9797 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15249), .ZN(n15259) );
  XNOR2_X1 U9798 ( .A(n8650), .B(n7484), .ZN(n15258) );
  NOR2_X1 U9799 ( .A1(n15259), .A2(n15258), .ZN(n15257) );
  NAND2_X1 U9800 ( .A1(n14707), .A2(n14706), .ZN(n14705) );
  NAND2_X1 U9801 ( .A1(n15255), .A2(n15254), .ZN(n7486) );
  AOI21_X1 U9802 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n7486), .A(n15253), .ZN(
        n15245) );
  XNOR2_X1 U9803 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n7489), .ZN(n7491) );
  NAND2_X1 U9804 ( .A1(n7490), .A2(n7491), .ZN(n7492) );
  INV_X1 U9805 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15247) );
  INV_X1 U9806 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7493) );
  NOR2_X1 U9807 ( .A1(n7494), .A2(n7493), .ZN(n7497) );
  XNOR2_X1 U9808 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n7496) );
  XOR2_X1 U9809 ( .A(n7496), .B(n7495), .Z(n14710) );
  INV_X1 U9810 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7500) );
  XNOR2_X1 U9811 ( .A(n7498), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15252) );
  XNOR2_X1 U9812 ( .A(n7502), .B(n7501), .ZN(n7504) );
  NAND2_X1 U9813 ( .A1(n7503), .A2(n7504), .ZN(n7505) );
  INV_X1 U9814 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n15044) );
  NOR2_X1 U9815 ( .A1(n7506), .A2(n7507), .ZN(n7508) );
  INV_X1 U9816 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14716) );
  XNOR2_X1 U9817 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n7509), .ZN(n14718) );
  NAND2_X1 U9818 ( .A1(n14719), .A2(n14718), .ZN(n7510) );
  NOR2_X1 U9819 ( .A1(n14719), .A2(n14718), .ZN(n14717) );
  NAND2_X1 U9820 ( .A1(n14845), .A2(n14844), .ZN(n14843) );
  NAND2_X1 U9821 ( .A1(n14849), .A2(n14848), .ZN(n7511) );
  XNOR2_X1 U9822 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7513) );
  XOR2_X1 U9823 ( .A(n7513), .B(n7512), .Z(n14852) );
  XOR2_X1 U9824 ( .A(n7515), .B(n7514), .Z(n7517) );
  INV_X1 U9825 ( .A(n14856), .ZN(n14857) );
  INV_X1 U9826 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14859) );
  INV_X1 U9827 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14864) );
  INV_X1 U9828 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14753) );
  NAND2_X1 U9829 ( .A1(n7522), .A2(n7521), .ZN(n7523) );
  INV_X1 U9830 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n7527) );
  NAND2_X1 U9831 ( .A1(n7525), .A2(n7524), .ZN(n7526) );
  OAI21_X1 U9832 ( .B1(n7527), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n7526), .ZN(
        n7528) );
  XNOR2_X1 U9833 ( .A(n7528), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n7530) );
  XNOR2_X1 U9834 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7529) );
  XNOR2_X1 U9835 ( .A(n7530), .B(n7529), .ZN(n7531) );
  NAND2_X1 U9836 ( .A1(n8598), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7698) );
  INV_X1 U9837 ( .A(n7698), .ZN(n7533) );
  NAND2_X1 U9838 ( .A1(n7534), .A2(n7533), .ZN(n7700) );
  NAND2_X1 U9839 ( .A1(n8669), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7535) );
  NAND2_X1 U9840 ( .A1(n7700), .A2(n7535), .ZN(n7719) );
  NAND2_X1 U9841 ( .A1(n8846), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7537) );
  NAND2_X1 U9842 ( .A1(n13734), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7536) );
  AND2_X1 U9843 ( .A1(n7537), .A2(n7536), .ZN(n7718) );
  NAND2_X1 U9844 ( .A1(n7719), .A2(n7718), .ZN(n7538) );
  NAND2_X1 U9845 ( .A1(n8850), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7540) );
  INV_X1 U9846 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9219) );
  NAND2_X1 U9847 ( .A1(n9219), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7539) );
  NAND2_X1 U9848 ( .A1(n8246), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7542) );
  INV_X1 U9849 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n8296) );
  NAND2_X1 U9850 ( .A1(n8296), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7541) );
  NAND2_X1 U9851 ( .A1(n6771), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7545) );
  INV_X1 U9852 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n8334) );
  NAND2_X1 U9853 ( .A1(n8334), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7544) );
  NAND2_X1 U9854 ( .A1(n8308), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7546) );
  NAND2_X1 U9855 ( .A1(n13735), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7548) );
  NAND2_X1 U9856 ( .A1(n8318), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n7547) );
  NAND2_X1 U9857 ( .A1(n7548), .A2(n7547), .ZN(n7789) );
  NAND2_X1 U9858 ( .A1(n8365), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7551) );
  INV_X1 U9859 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7549) );
  NAND2_X1 U9860 ( .A1(n7549), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n7550) );
  NAND2_X1 U9861 ( .A1(n7814), .A2(n7551), .ZN(n7842) );
  NAND2_X1 U9862 ( .A1(n8377), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7553) );
  NAND2_X1 U9863 ( .A1(n8382), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n7552) );
  NAND2_X1 U9864 ( .A1(n7842), .A2(n7841), .ZN(n7844) );
  NAND2_X1 U9865 ( .A1(n7844), .A2(n7553), .ZN(n7825) );
  NAND2_X1 U9866 ( .A1(n8472), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7555) );
  NAND2_X1 U9867 ( .A1(n8469), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n7554) );
  NAND2_X1 U9868 ( .A1(n7825), .A2(n7824), .ZN(n7827) );
  NAND2_X1 U9869 ( .A1(n7827), .A2(n7555), .ZN(n7865) );
  NAND2_X1 U9870 ( .A1(n8640), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7557) );
  NAND2_X1 U9871 ( .A1(n8633), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7556) );
  NAND2_X1 U9872 ( .A1(n7865), .A2(n7864), .ZN(n7867) );
  NAND2_X1 U9873 ( .A1(n7867), .A2(n7557), .ZN(n7883) );
  NAND2_X1 U9874 ( .A1(n8835), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7559) );
  NAND2_X1 U9875 ( .A1(n8840), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7558) );
  NAND2_X1 U9876 ( .A1(n9083), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7564) );
  NAND2_X1 U9877 ( .A1(n9080), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7563) );
  NAND2_X1 U9878 ( .A1(n9428), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7566) );
  NAND2_X1 U9879 ( .A1(n9415), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7565) );
  NAND2_X1 U9880 ( .A1(n9541), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7568) );
  NAND2_X1 U9881 ( .A1(n13726), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n7567) );
  NAND2_X1 U9882 ( .A1(n9588), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7570) );
  INV_X1 U9883 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U9884 ( .A1(n9596), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7569) );
  NAND2_X1 U9885 ( .A1(n10087), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7572) );
  NAND2_X1 U9886 ( .A1(n10083), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n7571) );
  INV_X1 U9887 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10259) );
  NAND2_X1 U9888 ( .A1(n10259), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n7574) );
  INV_X1 U9889 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10202) );
  NAND2_X1 U9890 ( .A1(n10202), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n7573) );
  INV_X1 U9891 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n13655) );
  NAND2_X1 U9892 ( .A1(n13655), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7578) );
  INV_X1 U9893 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n13615) );
  NAND2_X1 U9894 ( .A1(n13615), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7577) );
  AND2_X1 U9895 ( .A1(n7578), .A2(n7577), .ZN(n7968) );
  INV_X1 U9896 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10746) );
  XNOR2_X1 U9897 ( .A(n10746), .B(P1_DATAO_REG_22__SCAN_IN), .ZN(n7641) );
  INV_X1 U9898 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11538) );
  XNOR2_X1 U9899 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .ZN(n7982) );
  NAND2_X1 U9900 ( .A1(n7983), .A2(n7982), .ZN(n7580) );
  INV_X1 U9901 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11551) );
  NAND2_X1 U9902 ( .A1(n11551), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7579) );
  NAND2_X1 U9903 ( .A1(n7581), .A2(n11565), .ZN(n7582) );
  INV_X1 U9904 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n14087) );
  NAND2_X1 U9905 ( .A1(n14087), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7584) );
  INV_X1 U9906 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7585) );
  NAND2_X1 U9907 ( .A1(n7585), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7586) );
  INV_X1 U9908 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14688) );
  AND2_X1 U9909 ( .A1(n14688), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7587) );
  INV_X1 U9910 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14083) );
  NAND2_X1 U9911 ( .A1(n14083), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7588) );
  XNOR2_X1 U9912 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n7589) );
  XNOR2_X1 U9913 ( .A(n11649), .B(n7589), .ZN(n12509) );
  NOR2_X2 U9914 ( .A1(n7878), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n7681) );
  NOR2_X1 U9915 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), .ZN(
        n7601) );
  INV_X1 U9916 ( .A(n7614), .ZN(n7604) );
  NAND2_X4 U9917 ( .A1(n8044), .A2(n8045), .ZN(n9135) );
  NAND2_X1 U9918 ( .A1(n12509), .A2(n12748), .ZN(n7609) );
  INV_X1 U9919 ( .A(SI_27_), .ZN(n12511) );
  OR2_X1 U9920 ( .A1(n6422), .A2(n12511), .ZN(n7608) );
  INV_X1 U9921 ( .A(n7618), .ZN(n12506) );
  INV_X1 U9922 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7613) );
  NAND2_X1 U9923 ( .A1(n7612), .A2(n7617), .ZN(n13397) );
  INV_X1 U9924 ( .A(n13397), .ZN(n7619) );
  AND2_X2 U9925 ( .A1(n12506), .A2(n7619), .ZN(n7974) );
  NAND2_X1 U9926 ( .A1(n9876), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n7635) );
  AND2_X2 U9927 ( .A1(n7618), .A2(n13397), .ZN(n7711) );
  NAND2_X1 U9928 ( .A1(n10035), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n7634) );
  AND2_X4 U9929 ( .A1(n7618), .A2(n7619), .ZN(n7856) );
  INV_X1 U9930 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n7621) );
  NOR2_X1 U9931 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7754) );
  NAND2_X1 U9932 ( .A1(n7754), .A2(n9379), .ZN(n7767) );
  NAND2_X1 U9933 ( .A1(n7831), .A2(n7830), .ZN(n7833) );
  NAND2_X1 U9934 ( .A1(n7872), .A2(n7686), .ZN(n7902) );
  NOR2_X2 U9935 ( .A1(n7917), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7934) );
  NAND2_X1 U9936 ( .A1(n12651), .A2(n7934), .ZN(n7950) );
  INV_X1 U9937 ( .A(n7950), .ZN(n7620) );
  NAND2_X1 U9938 ( .A1(n7621), .A2(n7620), .ZN(n7952) );
  INV_X1 U9939 ( .A(n7952), .ZN(n7623) );
  INV_X1 U9940 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n7622) );
  INV_X1 U9941 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n7624) );
  INV_X1 U9942 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n13689) );
  INV_X1 U9943 ( .A(n8008), .ZN(n7628) );
  INV_X1 U9944 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n7627) );
  NAND2_X1 U9945 ( .A1(n7628), .A2(n7627), .ZN(n8018) );
  INV_X1 U9946 ( .A(n8018), .ZN(n7630) );
  INV_X1 U9947 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n7629) );
  NAND2_X1 U9948 ( .A1(n7630), .A2(n7629), .ZN(n8020) );
  NAND2_X1 U9949 ( .A1(n8020), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n7631) );
  NAND2_X1 U9950 ( .A1(n8038), .A2(n7631), .ZN(n13099) );
  NAND2_X1 U9951 ( .A1(n7856), .A2(n13099), .ZN(n7633) );
  NAND2_X1 U9952 ( .A1(n7852), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n7632) );
  NAND2_X1 U9953 ( .A1(n10035), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n7640) );
  NAND2_X1 U9954 ( .A1(n7852), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n7639) );
  NAND2_X1 U9955 ( .A1(n7977), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n7636) );
  NAND2_X1 U9956 ( .A1(n7986), .A2(n7636), .ZN(n13167) );
  NAND2_X1 U9957 ( .A1(n7856), .A2(n13167), .ZN(n7638) );
  NAND2_X1 U9958 ( .A1(n7974), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n7637) );
  XNOR2_X1 U9959 ( .A(n7642), .B(n7641), .ZN(n9829) );
  NAND2_X1 U9960 ( .A1(n9829), .A2(n12748), .ZN(n7644) );
  NAND2_X1 U9961 ( .A1(n8005), .A2(SI_22_), .ZN(n7643) );
  NAND2_X1 U9962 ( .A1(n10035), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n7649) );
  NAND2_X1 U9963 ( .A1(n7852), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n7648) );
  NAND2_X1 U9964 ( .A1(n7673), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7645) );
  NAND2_X1 U9965 ( .A1(n7962), .A2(n7645), .ZN(n13203) );
  NAND2_X1 U9966 ( .A1(n7856), .A2(n13203), .ZN(n7647) );
  NAND2_X1 U9967 ( .A1(n7974), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n7646) );
  NAND4_X1 U9968 ( .A1(n7649), .A2(n7648), .A3(n7647), .A4(n7646), .ZN(n13184)
         );
  INV_X1 U9969 ( .A(n13184), .ZN(n13211) );
  OR2_X1 U9970 ( .A1(n7651), .A2(n7650), .ZN(n7652) );
  NAND2_X1 U9971 ( .A1(n7653), .A2(n7652), .ZN(n9017) );
  NAND2_X1 U9972 ( .A1(n9017), .A2(n12748), .ZN(n7663) );
  NAND2_X1 U9973 ( .A1(n7655), .A2(n7656), .ZN(n7913) );
  INV_X1 U9974 ( .A(n7913), .ZN(n7658) );
  NAND2_X1 U9975 ( .A1(n7658), .A2(n7657), .ZN(n7929) );
  AOI22_X1 U9976 ( .A1(n8005), .A2(n10198), .B1(n7947), .B2(n9776), .ZN(n7662)
         );
  OR2_X1 U9977 ( .A1(n7665), .A2(n7664), .ZN(n7666) );
  NAND2_X1 U9978 ( .A1(n7667), .A2(n7666), .ZN(n8826) );
  OR2_X1 U9979 ( .A1(n8826), .A2(n7749), .ZN(n7671) );
  NAND2_X1 U9980 ( .A1(n7668), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7669) );
  XNOR2_X1 U9981 ( .A(n7669), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13058) );
  AOI22_X1 U9982 ( .A1(n8005), .A2(SI_18_), .B1(n7947), .B2(n13058), .ZN(n7670) );
  NAND2_X1 U9983 ( .A1(n7671), .A2(n7670), .ZN(n12535) );
  INV_X1 U9984 ( .A(n12535), .ZN(n13371) );
  NAND2_X1 U9985 ( .A1(n9876), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n7677) );
  INV_X1 U9986 ( .A(n7711), .ZN(n7725) );
  INV_X1 U9987 ( .A(n7725), .ZN(n10035) );
  NAND2_X1 U9988 ( .A1(n10035), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7676) );
  NAND2_X1 U9989 ( .A1(n7952), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7672) );
  NAND2_X1 U9990 ( .A1(n7673), .A2(n7672), .ZN(n13215) );
  NAND2_X1 U9991 ( .A1(n7856), .A2(n13215), .ZN(n7675) );
  NAND2_X1 U9992 ( .A1(n7852), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n7674) );
  NAND4_X1 U9993 ( .A1(n7677), .A2(n7676), .A3(n7675), .A4(n7674), .ZN(n13222)
         );
  NAND2_X1 U9994 ( .A1(n7678), .A2(n9045), .ZN(n7679) );
  NAND2_X1 U9995 ( .A1(n7680), .A2(n7679), .ZN(n8383) );
  NAND2_X1 U9996 ( .A1(n8383), .A2(n12748), .ZN(n7685) );
  BUF_X1 U9997 ( .A(n7681), .Z(n7682) );
  INV_X1 U9998 ( .A(n7682), .ZN(n7880) );
  NAND2_X1 U9999 ( .A1(n7880), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7683) );
  XNOR2_X1 U10000 ( .A(n7683), .B(n7595), .ZN(n11127) );
  AOI22_X1 U10001 ( .A1(n8005), .A2(n9033), .B1(n7947), .B2(n11127), .ZN(n7684) );
  NAND2_X1 U10002 ( .A1(n7685), .A2(n7684), .ZN(n14755) );
  INV_X1 U10003 ( .A(n14755), .ZN(n13257) );
  OR2_X1 U10004 ( .A1(n7872), .A2(n7686), .ZN(n7687) );
  AND2_X1 U10005 ( .A1(n7687), .A2(n7902), .ZN(n14768) );
  INV_X1 U10006 ( .A(n14768), .ZN(n12684) );
  NAND2_X1 U10007 ( .A1(n7856), .A2(n12684), .ZN(n7691) );
  NAND2_X1 U10008 ( .A1(n7711), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7690) );
  NAND2_X1 U10009 ( .A1(n7852), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7689) );
  NAND2_X1 U10010 ( .A1(n9876), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7688) );
  NAND4_X1 U10011 ( .A1(n7691), .A2(n7690), .A3(n7689), .A4(n7688), .ZN(n13262) );
  NAND2_X1 U10012 ( .A1(n7852), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7695) );
  NAND2_X1 U10013 ( .A1(n7974), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7694) );
  NAND2_X1 U10014 ( .A1(n7711), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7693) );
  NAND2_X1 U10015 ( .A1(n7856), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7692) );
  INV_X1 U10016 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7697) );
  NAND2_X1 U10017 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n7696) );
  XNOR2_X1 U10018 ( .A(n7697), .B(n7696), .ZN(n9173) );
  NAND2_X1 U10019 ( .A1(n7699), .A2(n7698), .ZN(n7701) );
  AND2_X1 U10020 ( .A1(n7701), .A2(n7700), .ZN(n8267) );
  NAND2_X1 U10021 ( .A1(n9780), .A2(n9779), .ZN(n12775) );
  NAND2_X1 U10022 ( .A1(n7711), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7706) );
  NAND2_X1 U10023 ( .A1(n7852), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7705) );
  NAND2_X1 U10024 ( .A1(n7974), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7704) );
  NAND2_X1 U10025 ( .A1(n7856), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7703) );
  NAND4_X2 U10026 ( .A1(n7706), .A2(n7705), .A3(n7704), .A4(n7703), .ZN(n15193) );
  INV_X1 U10027 ( .A(SI_0_), .ZN(n8705) );
  OR2_X1 U10028 ( .A1(n7750), .A2(n8705), .ZN(n7709) );
  XNOR2_X1 U10029 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(P2_DATAO_REG_0__SCAN_IN), 
        .ZN(n8273) );
  NAND2_X1 U10030 ( .A1(n7947), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n7707) );
  INV_X1 U10031 ( .A(n12771), .ZN(n9675) );
  NAND2_X1 U10032 ( .A1(n15193), .A2(n9675), .ZN(n15188) );
  INV_X1 U10033 ( .A(n15188), .ZN(n9822) );
  NAND2_X1 U10034 ( .A1(n9780), .A2(n15187), .ZN(n7710) );
  NAND2_X1 U10035 ( .A1(n7856), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7715) );
  NAND2_X1 U10036 ( .A1(n7711), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7714) );
  NAND2_X1 U10037 ( .A1(n7974), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7712) );
  OR2_X1 U10038 ( .A1(n7716), .A2(n7613), .ZN(n7717) );
  XNOR2_X1 U10039 ( .A(n7719), .B(n7718), .ZN(n8202) );
  OR2_X1 U10040 ( .A1(n7749), .A2(n8202), .ZN(n7721) );
  OR2_X1 U10041 ( .A1(n6422), .A2(SI_2_), .ZN(n7720) );
  OAI211_X1 U10042 ( .C1(n9207), .C2(n9135), .A(n7721), .B(n7720), .ZN(n7722)
         );
  INV_X1 U10043 ( .A(n7722), .ZN(n9778) );
  NAND2_X1 U10044 ( .A1(n15194), .A2(n7722), .ZN(n12778) );
  AND2_X2 U10045 ( .A1(n12777), .A2(n12778), .ZN(n15175) );
  INV_X1 U10046 ( .A(n15175), .ZN(n12774) );
  NOR2_X1 U10047 ( .A1(n15194), .A2(n9778), .ZN(n7723) );
  AOI21_X1 U10048 ( .B1(n15171), .B2(n12774), .A(n7723), .ZN(n10048) );
  INV_X1 U10049 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n7724) );
  NAND2_X1 U10050 ( .A1(n7856), .A2(n7724), .ZN(n7729) );
  NAND2_X1 U10051 ( .A1(n7711), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7728) );
  NAND2_X1 U10052 ( .A1(n7852), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7727) );
  NAND2_X1 U10053 ( .A1(n7974), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7726) );
  NAND4_X1 U10054 ( .A1(n7729), .A2(n7728), .A3(n7727), .A4(n7726), .ZN(n15172) );
  NAND2_X1 U10055 ( .A1(n7730), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7731) );
  XNOR2_X1 U10056 ( .A(n7731), .B(P3_IR_REG_3__SCAN_IN), .ZN(n9478) );
  XNOR2_X1 U10057 ( .A(n7733), .B(n7732), .ZN(n8196) );
  OR2_X1 U10058 ( .A1(n7749), .A2(n8196), .ZN(n7735) );
  OR2_X1 U10059 ( .A1(n6422), .A2(SI_3_), .ZN(n7734) );
  OAI211_X1 U10060 ( .C1(n9478), .C2(n9135), .A(n7735), .B(n7734), .ZN(n10495)
         );
  INV_X1 U10061 ( .A(n10495), .ZN(n10052) );
  NAND2_X1 U10062 ( .A1(n10093), .A2(n10052), .ZN(n12785) );
  NAND2_X1 U10063 ( .A1(n15172), .A2(n10495), .ZN(n12784) );
  AND2_X1 U10064 ( .A1(n12785), .A2(n12784), .ZN(n12929) );
  INV_X1 U10065 ( .A(n12929), .ZN(n10047) );
  NAND2_X1 U10066 ( .A1(n10048), .A2(n10047), .ZN(n10046) );
  NAND2_X1 U10067 ( .A1(n15172), .A2(n10052), .ZN(n7736) );
  NAND2_X1 U10068 ( .A1(n10046), .A2(n7736), .ZN(n10146) );
  NAND2_X1 U10069 ( .A1(n9876), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7741) );
  NAND2_X1 U10070 ( .A1(n7711), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7740) );
  AND2_X1 U10071 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7737) );
  OR2_X1 U10072 ( .A1(n7737), .A2(n7754), .ZN(n10088) );
  NAND2_X1 U10073 ( .A1(n7856), .A2(n10088), .ZN(n7739) );
  NAND2_X1 U10074 ( .A1(n7852), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7738) );
  NAND4_X1 U10075 ( .A1(n7741), .A2(n7740), .A3(n7739), .A4(n7738), .ZN(n12975) );
  NAND2_X1 U10076 ( .A1(n7742), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7743) );
  MUX2_X1 U10077 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7743), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n7746) );
  INV_X1 U10078 ( .A(n7744), .ZN(n7745) );
  XNOR2_X1 U10079 ( .A(n7748), .B(n7747), .ZN(n8188) );
  OR2_X1 U10080 ( .A1(n7749), .A2(n8188), .ZN(n7752) );
  OR2_X1 U10081 ( .A1(n6422), .A2(SI_4_), .ZN(n7751) );
  OAI211_X1 U10082 ( .C1(n9190), .C2(n9135), .A(n7752), .B(n7751), .ZN(n12787)
         );
  INV_X1 U10083 ( .A(n12787), .ZN(n10491) );
  XNOR2_X1 U10084 ( .A(n12975), .B(n10491), .ZN(n12937) );
  INV_X1 U10085 ( .A(n12937), .ZN(n10145) );
  NAND2_X1 U10086 ( .A1(n10146), .A2(n10145), .ZN(n10144) );
  NAND2_X1 U10087 ( .A1(n12975), .A2(n10491), .ZN(n7753) );
  NAND2_X1 U10088 ( .A1(n10144), .A2(n7753), .ZN(n10576) );
  NAND2_X1 U10089 ( .A1(n9876), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7759) );
  NAND2_X1 U10090 ( .A1(n7711), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7758) );
  OR2_X1 U10091 ( .A1(n7754), .A2(n9379), .ZN(n7755) );
  NAND2_X1 U10092 ( .A1(n7767), .A2(n7755), .ZN(n10584) );
  NAND2_X1 U10093 ( .A1(n7856), .A2(n10584), .ZN(n7757) );
  NAND2_X1 U10094 ( .A1(n7852), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7756) );
  NAND4_X1 U10095 ( .A1(n7759), .A2(n7758), .A3(n7757), .A4(n7756), .ZN(n12974) );
  INV_X1 U10096 ( .A(n12974), .ZN(n7766) );
  OR2_X1 U10097 ( .A1(n7744), .A2(n7613), .ZN(n7760) );
  XNOR2_X1 U10098 ( .A(n7760), .B(P3_IR_REG_5__SCAN_IN), .ZN(n9384) );
  XNOR2_X1 U10099 ( .A(n7762), .B(n7761), .ZN(n8191) );
  OR2_X1 U10100 ( .A1(n7749), .A2(n8191), .ZN(n7764) );
  OR2_X1 U10101 ( .A1(n6422), .A2(SI_5_), .ZN(n7763) );
  OAI211_X1 U10102 ( .C1(n9384), .C2(n9135), .A(n7764), .B(n7763), .ZN(n10583)
         );
  INV_X1 U10103 ( .A(n10583), .ZN(n7765) );
  NAND2_X1 U10104 ( .A1(n7766), .A2(n7765), .ZN(n12793) );
  NAND2_X1 U10105 ( .A1(n12974), .A2(n10583), .ZN(n12798) );
  NAND2_X1 U10106 ( .A1(n7766), .A2(n10583), .ZN(n10449) );
  NAND2_X1 U10107 ( .A1(n9876), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7772) );
  NAND2_X1 U10108 ( .A1(n7711), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7771) );
  NAND2_X1 U10109 ( .A1(n7767), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7768) );
  NAND2_X1 U10110 ( .A1(n7780), .A2(n7768), .ZN(n10677) );
  NAND2_X1 U10111 ( .A1(n7856), .A2(n10677), .ZN(n7770) );
  NAND2_X1 U10112 ( .A1(n7852), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7769) );
  NAND4_X1 U10113 ( .A1(n7772), .A2(n7771), .A3(n7770), .A4(n7769), .ZN(n12973) );
  INV_X1 U10114 ( .A(n12973), .ZN(n10618) );
  OR2_X1 U10115 ( .A1(n7773), .A2(n7613), .ZN(n7774) );
  XNOR2_X1 U10116 ( .A(n7774), .B(n7786), .ZN(n15127) );
  INV_X1 U10117 ( .A(SI_6_), .ZN(n8194) );
  OR2_X1 U10118 ( .A1(n6422), .A2(n8194), .ZN(n7778) );
  XNOR2_X1 U10119 ( .A(n8308), .B(P1_DATAO_REG_6__SCAN_IN), .ZN(n7775) );
  XNOR2_X1 U10120 ( .A(n7776), .B(n7775), .ZN(n8195) );
  OR2_X1 U10121 ( .A1(n7749), .A2(n8195), .ZN(n7777) );
  OAI211_X1 U10122 ( .C1(n9135), .C2(n15127), .A(n7778), .B(n7777), .ZN(n10669) );
  NAND2_X1 U10123 ( .A1(n10618), .A2(n10669), .ZN(n12800) );
  INV_X1 U10124 ( .A(n10669), .ZN(n10642) );
  NAND2_X1 U10125 ( .A1(n12973), .A2(n10642), .ZN(n12799) );
  INV_X1 U10126 ( .A(n12928), .ZN(n7779) );
  AND2_X1 U10127 ( .A1(n10449), .A2(n7779), .ZN(n10448) );
  NAND2_X1 U10128 ( .A1(n9876), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7785) );
  NAND2_X1 U10129 ( .A1(n10035), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7784) );
  AND2_X1 U10130 ( .A1(n7780), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7781) );
  OR2_X1 U10131 ( .A1(n7781), .A2(n7800), .ZN(n10609) );
  NAND2_X1 U10132 ( .A1(n7856), .A2(n10609), .ZN(n7783) );
  NAND2_X1 U10133 ( .A1(n7852), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7782) );
  NAND4_X1 U10134 ( .A1(n7785), .A2(n7784), .A3(n7783), .A4(n7782), .ZN(n12972) );
  NAND2_X1 U10135 ( .A1(n7773), .A2(n7786), .ZN(n7806) );
  NAND2_X1 U10136 ( .A1(n7806), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7788) );
  XNOR2_X1 U10137 ( .A(n7788), .B(n7787), .ZN(n10164) );
  INV_X1 U10138 ( .A(n10164), .ZN(n9984) );
  NAND2_X1 U10139 ( .A1(n7790), .A2(n7789), .ZN(n7791) );
  AND2_X1 U10140 ( .A1(n7792), .A2(n7791), .ZN(n8199) );
  OR2_X1 U10141 ( .A1(n7749), .A2(n8199), .ZN(n7794) );
  OR2_X1 U10142 ( .A1(n6422), .A2(SI_7_), .ZN(n7793) );
  OAI211_X1 U10143 ( .C1(n9984), .C2(n9135), .A(n7794), .B(n7793), .ZN(n12806)
         );
  XNOR2_X1 U10144 ( .A(n12972), .B(n12806), .ZN(n12933) );
  AND2_X1 U10145 ( .A1(n10448), .A2(n12933), .ZN(n7798) );
  INV_X1 U10146 ( .A(n12933), .ZN(n7795) );
  NAND2_X1 U10147 ( .A1(n12973), .A2(n10669), .ZN(n10598) );
  OR2_X1 U10148 ( .A1(n7795), .A2(n10598), .ZN(n7796) );
  NAND2_X1 U10149 ( .A1(n9876), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7805) );
  NAND2_X1 U10150 ( .A1(n10035), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7804) );
  NOR2_X1 U10151 ( .A1(n7800), .A2(n7799), .ZN(n7801) );
  OR2_X1 U10152 ( .A1(n7831), .A2(n7801), .ZN(n10823) );
  NAND2_X1 U10153 ( .A1(n7856), .A2(n10823), .ZN(n7803) );
  NAND2_X1 U10154 ( .A1(n7852), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7802) );
  NAND4_X1 U10155 ( .A1(n7805), .A2(n7804), .A3(n7803), .A4(n7802), .ZN(n12971) );
  INV_X1 U10156 ( .A(n12971), .ZN(n10960) );
  NAND2_X1 U10157 ( .A1(n7809), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7808) );
  MUX2_X1 U10158 ( .A(n7808), .B(P3_IR_REG_31__SCAN_IN), .S(n7807), .Z(n7810)
         );
  NAND2_X1 U10159 ( .A1(n7810), .A2(n7838), .ZN(n15149) );
  INV_X1 U10160 ( .A(SI_8_), .ZN(n8271) );
  OR2_X1 U10161 ( .A1(n6422), .A2(n8271), .ZN(n7816) );
  OR2_X1 U10162 ( .A1(n7812), .A2(n7811), .ZN(n7813) );
  NAND2_X1 U10163 ( .A1(n7814), .A2(n7813), .ZN(n8272) );
  OR2_X1 U10164 ( .A1(n7749), .A2(n8272), .ZN(n7815) );
  OAI211_X1 U10165 ( .C1(n9135), .C2(n15149), .A(n7816), .B(n7815), .ZN(n10732) );
  NAND2_X1 U10166 ( .A1(n10960), .A2(n10732), .ZN(n12812) );
  INV_X1 U10167 ( .A(n10732), .ZN(n10822) );
  NAND2_X1 U10168 ( .A1(n12971), .A2(n10822), .ZN(n12811) );
  INV_X1 U10169 ( .A(n12806), .ZN(n8050) );
  NAND2_X1 U10170 ( .A1(n12972), .A2(n8050), .ZN(n10813) );
  AND2_X1 U10171 ( .A1(n10812), .A2(n10813), .ZN(n7888) );
  NAND2_X1 U10172 ( .A1(n9876), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7821) );
  NAND2_X1 U10173 ( .A1(n7711), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7820) );
  NAND2_X1 U10174 ( .A1(n7833), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7817) );
  NAND2_X1 U10175 ( .A1(n7853), .A2(n7817), .ZN(n12597) );
  NAND2_X1 U10176 ( .A1(n7856), .A2(n12597), .ZN(n7819) );
  NAND2_X1 U10177 ( .A1(n7852), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7818) );
  NAND4_X1 U10178 ( .A1(n7821), .A2(n7820), .A3(n7819), .A4(n7818), .ZN(n12969) );
  INV_X1 U10179 ( .A(n7838), .ZN(n7822) );
  INV_X1 U10180 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7839) );
  NAND2_X1 U10181 ( .A1(n7822), .A2(n7839), .ZN(n7861) );
  NAND2_X1 U10182 ( .A1(n7861), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7823) );
  XNOR2_X1 U10183 ( .A(n7823), .B(P3_IR_REG_10__SCAN_IN), .ZN(n10346) );
  OR2_X1 U10184 ( .A1(n6422), .A2(SI_10_), .ZN(n7829) );
  OR2_X1 U10185 ( .A1(n7825), .A2(n7824), .ZN(n7826) );
  AND2_X1 U10186 ( .A1(n7827), .A2(n7826), .ZN(n8287) );
  OR2_X1 U10187 ( .A1(n7749), .A2(n8287), .ZN(n7828) );
  OAI211_X1 U10188 ( .C1(n10346), .C2(n9135), .A(n7829), .B(n7828), .ZN(n15227) );
  INV_X1 U10189 ( .A(n15227), .ZN(n12588) );
  NAND2_X1 U10190 ( .A1(n12969), .A2(n12588), .ZN(n7848) );
  INV_X1 U10191 ( .A(n12969), .ZN(n14777) );
  NAND2_X1 U10192 ( .A1(n14777), .A2(n12588), .ZN(n12820) );
  NAND2_X1 U10193 ( .A1(n12969), .A2(n15227), .ZN(n12819) );
  NAND2_X1 U10194 ( .A1(n12820), .A2(n12819), .ZN(n10886) );
  INV_X1 U10195 ( .A(n10886), .ZN(n12927) );
  OR2_X1 U10196 ( .A1(n7831), .A2(n7830), .ZN(n7832) );
  AND2_X1 U10197 ( .A1(n7833), .A2(n7832), .ZN(n15170) );
  INV_X1 U10198 ( .A(n15170), .ZN(n10963) );
  NAND2_X1 U10199 ( .A1(n7856), .A2(n10963), .ZN(n7837) );
  NAND2_X1 U10200 ( .A1(n10035), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7836) );
  NAND2_X1 U10201 ( .A1(n7852), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7835) );
  NAND2_X1 U10202 ( .A1(n9876), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7834) );
  NAND4_X1 U10203 ( .A1(n7837), .A2(n7836), .A3(n7835), .A4(n7834), .ZN(n12970) );
  NAND2_X1 U10204 ( .A1(n7838), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7840) );
  XNOR2_X1 U10205 ( .A(n7840), .B(n7839), .ZN(n10343) );
  INV_X1 U10206 ( .A(n10343), .ZN(n7847) );
  OR2_X1 U10207 ( .A1(n6422), .A2(SI_9_), .ZN(n7846) );
  OR2_X1 U10208 ( .A1(n7842), .A2(n7841), .ZN(n7843) );
  AND2_X1 U10209 ( .A1(n7844), .A2(n7843), .ZN(n8268) );
  OR2_X1 U10210 ( .A1(n7749), .A2(n8268), .ZN(n7845) );
  OAI211_X1 U10211 ( .C1(n7847), .C2(n9135), .A(n7846), .B(n7845), .ZN(n15164)
         );
  INV_X1 U10212 ( .A(n15164), .ZN(n8052) );
  NAND2_X1 U10213 ( .A1(n12970), .A2(n8052), .ZN(n10882) );
  OR2_X1 U10214 ( .A1(n12927), .A2(n10882), .ZN(n10883) );
  AND2_X1 U10215 ( .A1(n7848), .A2(n10883), .ZN(n7891) );
  AND2_X1 U10216 ( .A1(n7888), .A2(n7891), .ZN(n7851) );
  INV_X1 U10217 ( .A(n7891), .ZN(n7850) );
  XNOR2_X1 U10218 ( .A(n12970), .B(n8052), .ZN(n12936) );
  INV_X1 U10219 ( .A(n12936), .ZN(n10992) );
  AND2_X1 U10220 ( .A1(n10992), .A2(n10886), .ZN(n7890) );
  NAND2_X1 U10221 ( .A1(n10960), .A2(n10822), .ZN(n7889) );
  AND2_X1 U10222 ( .A1(n7890), .A2(n7889), .ZN(n7849) );
  AOI21_X1 U10223 ( .B1(n10814), .B2(n7851), .A(n7402), .ZN(n7870) );
  NAND2_X1 U10224 ( .A1(n7711), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7860) );
  NAND2_X1 U10225 ( .A1(n7852), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7859) );
  NAND2_X1 U10226 ( .A1(n9876), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7858) );
  NAND2_X1 U10227 ( .A1(n7853), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7854) );
  AND2_X1 U10228 ( .A1(n7871), .A2(n7854), .ZN(n14783) );
  INV_X1 U10229 ( .A(n14783), .ZN(n7855) );
  NAND2_X1 U10230 ( .A1(n7856), .A2(n7855), .ZN(n7857) );
  NAND4_X1 U10231 ( .A1(n7860), .A2(n7859), .A3(n7858), .A4(n7857), .ZN(n12968) );
  OAI21_X1 U10232 ( .B1(n7861), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7863) );
  INV_X1 U10233 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7862) );
  XNOR2_X1 U10234 ( .A(n7863), .B(n7862), .ZN(n10789) );
  OR2_X1 U10235 ( .A1(n6422), .A2(SI_11_), .ZN(n7869) );
  OR2_X1 U10236 ( .A1(n7865), .A2(n7864), .ZN(n7866) );
  AND2_X1 U10237 ( .A1(n7867), .A2(n7866), .ZN(n8314) );
  OR2_X1 U10238 ( .A1(n7749), .A2(n8314), .ZN(n7868) );
  OAI211_X1 U10239 ( .C1(n10767), .C2(n9135), .A(n7869), .B(n7868), .ZN(n14769) );
  INV_X1 U10240 ( .A(n14769), .ZN(n8057) );
  OAI21_X1 U10241 ( .B1(n7870), .B2(n12968), .A(n8057), .ZN(n11094) );
  AND2_X1 U10242 ( .A1(n7871), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7873) );
  OR2_X1 U10243 ( .A1(n7873), .A2(n7872), .ZN(n12637) );
  NAND2_X1 U10244 ( .A1(n7856), .A2(n12637), .ZN(n7877) );
  NAND2_X1 U10245 ( .A1(n10035), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7876) );
  NAND2_X1 U10246 ( .A1(n7852), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7875) );
  NAND2_X1 U10247 ( .A1(n9876), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7874) );
  NAND2_X1 U10248 ( .A1(n7878), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7879) );
  MUX2_X1 U10249 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7879), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n7881) );
  NAND2_X1 U10250 ( .A1(n7881), .A2(n7880), .ZN(n12985) );
  OR2_X1 U10251 ( .A1(n7883), .A2(n7882), .ZN(n7884) );
  NAND2_X1 U10252 ( .A1(n7885), .A2(n7884), .ZN(n8362) );
  OR2_X1 U10253 ( .A1(n8362), .A2(n7749), .ZN(n7887) );
  NAND2_X1 U10254 ( .A1(n8005), .A2(SI_12_), .ZN(n7886) );
  OAI211_X1 U10255 ( .C1(n9135), .C2(n12985), .A(n7887), .B(n7886), .ZN(n12634) );
  INV_X1 U10256 ( .A(n12634), .ZN(n14789) );
  OR2_X1 U10257 ( .A1(n14775), .A2(n14789), .ZN(n7892) );
  AND2_X1 U10258 ( .A1(n11094), .A2(n7892), .ZN(n7894) );
  NAND2_X1 U10259 ( .A1(n10884), .A2(n7891), .ZN(n14773) );
  NAND2_X1 U10260 ( .A1(n14773), .A2(n12968), .ZN(n11095) );
  INV_X1 U10261 ( .A(n7892), .ZN(n7893) );
  OR2_X1 U10262 ( .A1(n14775), .A2(n12634), .ZN(n12830) );
  NAND2_X1 U10263 ( .A1(n14775), .A2(n12634), .ZN(n12831) );
  OR2_X1 U10264 ( .A1(n7896), .A2(n7895), .ZN(n7897) );
  NAND2_X1 U10265 ( .A1(n7898), .A2(n7897), .ZN(n8443) );
  OR2_X1 U10266 ( .A1(n8443), .A2(n7749), .ZN(n7901) );
  OR2_X1 U10267 ( .A1(n7655), .A2(n7613), .ZN(n7899) );
  XNOR2_X1 U10268 ( .A(n7899), .B(P3_IR_REG_14__SCAN_IN), .ZN(n11122) );
  AOI22_X1 U10269 ( .A1(n8005), .A2(SI_14_), .B1(n7947), .B2(n11122), .ZN(
        n7900) );
  NAND2_X1 U10270 ( .A1(n7901), .A2(n7900), .ZN(n12579) );
  NAND2_X1 U10271 ( .A1(n9876), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7907) );
  NAND2_X1 U10272 ( .A1(n10035), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7906) );
  NAND2_X1 U10273 ( .A1(n7902), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7903) );
  NAND2_X1 U10274 ( .A1(n7917), .A2(n7903), .ZN(n13267) );
  NAND2_X1 U10275 ( .A1(n7856), .A2(n13267), .ZN(n7905) );
  NAND2_X1 U10276 ( .A1(n7852), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n7904) );
  NAND4_X1 U10277 ( .A1(n7907), .A2(n7906), .A3(n7905), .A4(n7904), .ZN(n14759) );
  OR2_X1 U10278 ( .A1(n12579), .A2(n13247), .ZN(n12844) );
  NAND2_X1 U10279 ( .A1(n12579), .A2(n13247), .ZN(n12843) );
  NAND3_X1 U10280 ( .A1(n13260), .A2(n13257), .A3(n13262), .ZN(n7908) );
  INV_X1 U10281 ( .A(n12579), .ZN(n13385) );
  OR2_X1 U10282 ( .A1(n7910), .A2(n7909), .ZN(n7911) );
  NAND2_X1 U10283 ( .A1(n7912), .A2(n7911), .ZN(n8560) );
  OR2_X1 U10284 ( .A1(n8560), .A2(n7749), .ZN(n7916) );
  NAND2_X1 U10285 ( .A1(n7913), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7914) );
  XNOR2_X1 U10286 ( .A(n7914), .B(P3_IR_REG_15__SCAN_IN), .ZN(n11272) );
  AOI22_X1 U10287 ( .A1(n8005), .A2(SI_15_), .B1(n7947), .B2(n11272), .ZN(
        n7915) );
  NAND2_X1 U10288 ( .A1(n7916), .A2(n7915), .ZN(n12736) );
  NAND2_X1 U10289 ( .A1(n9876), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7922) );
  NAND2_X1 U10290 ( .A1(n10035), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7921) );
  AND2_X1 U10291 ( .A1(n7917), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7918) );
  OR2_X1 U10292 ( .A1(n7918), .A2(n7934), .ZN(n13251) );
  NAND2_X1 U10293 ( .A1(n7856), .A2(n13251), .ZN(n7920) );
  NAND2_X1 U10294 ( .A1(n7852), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n7919) );
  INV_X1 U10295 ( .A(n12736), .ZN(n13380) );
  OR2_X1 U10296 ( .A1(n7926), .A2(n7925), .ZN(n7927) );
  NAND2_X1 U10297 ( .A1(n7928), .A2(n7927), .ZN(n8634) );
  OR2_X1 U10298 ( .A1(n8634), .A2(n7749), .ZN(n7933) );
  NAND2_X1 U10299 ( .A1(n7929), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7930) );
  MUX2_X1 U10300 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7930), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n7931) );
  AND2_X1 U10301 ( .A1(n7931), .A2(n7944), .ZN(n13018) );
  AOI22_X1 U10302 ( .A1(n8005), .A2(SI_16_), .B1(n7947), .B2(n13018), .ZN(
        n7932) );
  NAND2_X1 U10303 ( .A1(n7933), .A2(n7932), .ZN(n13239) );
  NAND2_X1 U10304 ( .A1(n9876), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7939) );
  NAND2_X1 U10305 ( .A1(n10035), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7938) );
  OR2_X1 U10306 ( .A1(n7934), .A2(n12651), .ZN(n7935) );
  NAND2_X1 U10307 ( .A1(n7935), .A2(n7950), .ZN(n13240) );
  NAND2_X1 U10308 ( .A1(n7856), .A2(n13240), .ZN(n7937) );
  NAND2_X1 U10309 ( .A1(n7852), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n7936) );
  NAND4_X1 U10310 ( .A1(n7939), .A2(n7938), .A3(n7937), .A4(n7936), .ZN(n13221) );
  OR2_X1 U10311 ( .A1(n13239), .A2(n13248), .ZN(n12854) );
  NAND2_X1 U10312 ( .A1(n13239), .A2(n13248), .ZN(n12853) );
  INV_X1 U10313 ( .A(n13237), .ZN(n13231) );
  OR2_X1 U10314 ( .A1(n7941), .A2(n7940), .ZN(n7942) );
  NAND2_X1 U10315 ( .A1(n7943), .A2(n7942), .ZN(n8759) );
  NAND2_X1 U10316 ( .A1(n8759), .A2(n12748), .ZN(n7949) );
  NAND2_X1 U10317 ( .A1(n7944), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7946) );
  AOI22_X1 U10318 ( .A1(n8005), .A2(n10080), .B1(n7947), .B2(n13044), .ZN(
        n7948) );
  NAND2_X1 U10319 ( .A1(n7949), .A2(n7948), .ZN(n13322) );
  NAND2_X1 U10320 ( .A1(n9876), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n7956) );
  NAND2_X1 U10321 ( .A1(n7711), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7955) );
  NAND2_X1 U10322 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(n7950), .ZN(n7951) );
  NAND2_X1 U10323 ( .A1(n7952), .A2(n7951), .ZN(n13227) );
  NAND2_X1 U10324 ( .A1(n7856), .A2(n13227), .ZN(n7954) );
  NAND2_X1 U10325 ( .A1(n7852), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n7953) );
  NAND4_X1 U10326 ( .A1(n7956), .A2(n7955), .A3(n7954), .A4(n7953), .ZN(n12966) );
  OR2_X1 U10327 ( .A1(n13322), .A2(n12966), .ZN(n12857) );
  NAND2_X1 U10328 ( .A1(n13322), .A2(n12966), .ZN(n12860) );
  INV_X1 U10329 ( .A(n12966), .ZN(n13234) );
  NAND2_X1 U10330 ( .A1(n12535), .A2(n12538), .ZN(n12863) );
  NAND2_X1 U10331 ( .A1(n12858), .A2(n12863), .ZN(n13214) );
  INV_X1 U10332 ( .A(n13214), .ZN(n13209) );
  NOR2_X1 U10333 ( .A1(n13309), .A2(n13184), .ZN(n8060) );
  INV_X1 U10334 ( .A(n8060), .ZN(n12868) );
  NAND2_X1 U10335 ( .A1(n13309), .A2(n13184), .ZN(n12869) );
  NAND2_X1 U10336 ( .A1(n12868), .A2(n12869), .ZN(n13198) );
  NAND2_X1 U10337 ( .A1(n13199), .A2(n13198), .ZN(n13197) );
  OAI21_X1 U10338 ( .B1(n13211), .B2(n13309), .A(n13197), .ZN(n13183) );
  NAND2_X1 U10339 ( .A1(n7957), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7958) );
  NAND2_X1 U10340 ( .A1(n7959), .A2(n7958), .ZN(n9501) );
  OR2_X1 U10341 ( .A1(n9501), .A2(n7749), .ZN(n7961) );
  INV_X1 U10342 ( .A(SI_20_), .ZN(n10185) );
  OR2_X1 U10343 ( .A1(n6422), .A2(n10185), .ZN(n7960) );
  NAND2_X2 U10344 ( .A1(n7961), .A2(n7960), .ZN(n13305) );
  NAND2_X1 U10345 ( .A1(n10035), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n7967) );
  NAND2_X1 U10346 ( .A1(n7974), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n7966) );
  NAND2_X1 U10347 ( .A1(n7962), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n7963) );
  NAND2_X1 U10348 ( .A1(n7975), .A2(n7963), .ZN(n13190) );
  NAND2_X1 U10349 ( .A1(n7856), .A2(n13190), .ZN(n7965) );
  NAND2_X1 U10350 ( .A1(n7852), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n7964) );
  NAND4_X1 U10351 ( .A1(n7967), .A2(n7966), .A3(n7965), .A4(n7964), .ZN(n13200) );
  NAND2_X1 U10352 ( .A1(n13305), .A2(n13174), .ZN(n12874) );
  INV_X1 U10353 ( .A(n13188), .ZN(n12944) );
  OR2_X1 U10354 ( .A1(n7969), .A2(n7968), .ZN(n7970) );
  NAND2_X1 U10355 ( .A1(n7971), .A2(n7970), .ZN(n9581) );
  OR2_X1 U10356 ( .A1(n9581), .A2(n7749), .ZN(n7973) );
  NAND2_X1 U10357 ( .A1(n8005), .A2(SI_21_), .ZN(n7972) );
  NAND2_X1 U10358 ( .A1(n7974), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n7981) );
  NAND2_X1 U10359 ( .A1(n7711), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n7980) );
  NAND2_X1 U10360 ( .A1(n7975), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n7976) );
  NAND2_X1 U10361 ( .A1(n7977), .A2(n7976), .ZN(n13178) );
  NAND2_X1 U10362 ( .A1(n7856), .A2(n13178), .ZN(n7979) );
  NAND2_X1 U10363 ( .A1(n7852), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n7978) );
  NAND4_X1 U10364 ( .A1(n7981), .A2(n7980), .A3(n7979), .A4(n7978), .ZN(n13185) );
  XNOR2_X1 U10365 ( .A(n7983), .B(n7982), .ZN(n10072) );
  NAND2_X1 U10366 ( .A1(n10072), .A2(n12748), .ZN(n7985) );
  INV_X1 U10367 ( .A(SI_23_), .ZN(n10074) );
  OR2_X1 U10368 ( .A1(n6422), .A2(n10074), .ZN(n7984) );
  NAND2_X1 U10369 ( .A1(n9876), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n7991) );
  NAND2_X1 U10370 ( .A1(n7711), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n7990) );
  NAND2_X1 U10371 ( .A1(n7986), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7987) );
  NAND2_X1 U10372 ( .A1(n7996), .A2(n7987), .ZN(n13156) );
  NAND2_X1 U10373 ( .A1(n7856), .A2(n13156), .ZN(n7989) );
  NAND2_X1 U10374 ( .A1(n7852), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n7988) );
  NAND2_X1 U10375 ( .A1(n13155), .A2(n13164), .ZN(n7992) );
  INV_X1 U10376 ( .A(n13148), .ZN(n7993) );
  AOI22_X2 U10377 ( .A1(n13149), .A2(n7993), .B1(n13136), .B2(n13155), .ZN(
        n13134) );
  INV_X1 U10378 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11163) );
  XNOR2_X1 U10379 ( .A(n7994), .B(n11163), .ZN(n11776) );
  NOR2_X1 U10380 ( .A1(n6422), .A2(n6925), .ZN(n7995) );
  AOI21_X2 U10381 ( .B1(n11776), .B2(n12748), .A(n7995), .ZN(n13289) );
  NAND2_X1 U10382 ( .A1(n9876), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8001) );
  NAND2_X1 U10383 ( .A1(n7711), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8000) );
  NAND2_X1 U10384 ( .A1(n7996), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n7997) );
  NAND2_X1 U10385 ( .A1(n8008), .A2(n7997), .ZN(n13141) );
  NAND2_X1 U10386 ( .A1(n7856), .A2(n13141), .ZN(n7999) );
  NAND2_X1 U10387 ( .A1(n7852), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n7998) );
  NAND4_X1 U10388 ( .A1(n8001), .A2(n8000), .A3(n7999), .A4(n7998), .ZN(n13151) );
  INV_X1 U10389 ( .A(n13151), .ZN(n12644) );
  NAND2_X1 U10390 ( .A1(n13289), .A2(n12644), .ZN(n8002) );
  XNOR2_X1 U10391 ( .A(n14087), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8003) );
  XNOR2_X1 U10392 ( .A(n8004), .B(n8003), .ZN(n10803) );
  NAND2_X1 U10393 ( .A1(n10803), .A2(n12748), .ZN(n8007) );
  NAND2_X1 U10394 ( .A1(n8005), .A2(SI_25_), .ZN(n8006) );
  NAND2_X1 U10395 ( .A1(n9876), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8013) );
  NAND2_X1 U10396 ( .A1(n7711), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8012) );
  NAND2_X1 U10397 ( .A1(n8008), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8009) );
  NAND2_X1 U10398 ( .A1(n8018), .A2(n8009), .ZN(n13129) );
  NAND2_X1 U10399 ( .A1(n7856), .A2(n13129), .ZN(n8011) );
  NAND2_X1 U10400 ( .A1(n7852), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8010) );
  NAND4_X1 U10401 ( .A1(n8013), .A2(n8012), .A3(n8011), .A4(n8010), .ZN(n13135) );
  NOR2_X1 U10402 ( .A1(n13128), .A2(n13110), .ZN(n8061) );
  INV_X1 U10403 ( .A(n8061), .ZN(n12889) );
  NAND2_X1 U10404 ( .A1(n13128), .A2(n13110), .ZN(n12890) );
  XNOR2_X1 U10405 ( .A(n14688), .B(P1_DATAO_REG_26__SCAN_IN), .ZN(n8014) );
  XNOR2_X1 U10406 ( .A(n8015), .B(n8014), .ZN(n10807) );
  NAND2_X1 U10407 ( .A1(n10807), .A2(n12748), .ZN(n8017) );
  INV_X1 U10408 ( .A(SI_26_), .ZN(n10810) );
  OR2_X1 U10409 ( .A1(n6422), .A2(n10810), .ZN(n8016) );
  NAND2_X1 U10410 ( .A1(n7711), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8024) );
  NAND2_X1 U10411 ( .A1(n7974), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8023) );
  NAND2_X1 U10412 ( .A1(n8018), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8019) );
  NAND2_X1 U10413 ( .A1(n8020), .A2(n8019), .ZN(n13117) );
  NAND2_X1 U10414 ( .A1(n7856), .A2(n13117), .ZN(n8022) );
  NAND2_X1 U10415 ( .A1(n7852), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8021) );
  NAND2_X1 U10416 ( .A1(n13348), .A2(n12565), .ZN(n8025) );
  NAND2_X1 U10417 ( .A1(n12564), .A2(n13125), .ZN(n8026) );
  INV_X1 U10418 ( .A(n11661), .ZN(n8027) );
  AOI21_X1 U10419 ( .B1(n12947), .B2(n8028), .A(n8027), .ZN(n8048) );
  NAND2_X1 U10420 ( .A1(n8068), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8031) );
  AND2_X1 U10421 ( .A1(n13072), .A2(n9830), .ZN(n8119) );
  NAND2_X1 U10422 ( .A1(n6469), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8032) );
  MUX2_X1 U10423 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8032), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8033) );
  AND2_X1 U10424 ( .A1(n8029), .A2(n8033), .ZN(n8117) );
  NAND2_X1 U10425 ( .A1(n8029), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8034) );
  MUX2_X1 U10426 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8034), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n8035) );
  NOR2_X1 U10427 ( .A1(n9775), .A2(n10042), .ZN(n12761) );
  NAND2_X1 U10428 ( .A1(n7974), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8043) );
  NAND2_X1 U10429 ( .A1(n7711), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8042) );
  INV_X1 U10430 ( .A(n8038), .ZN(n8037) );
  INV_X1 U10431 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8036) );
  NAND2_X1 U10432 ( .A1(n8037), .A2(n8036), .ZN(n11895) );
  NAND2_X1 U10433 ( .A1(n8038), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8039) );
  NAND2_X1 U10434 ( .A1(n11895), .A2(n8039), .ZN(n13093) );
  NAND2_X1 U10435 ( .A1(n7856), .A2(n13093), .ZN(n8041) );
  NAND2_X1 U10436 ( .A1(n7852), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8040) );
  INV_X1 U10437 ( .A(n12569), .ZN(n12965) );
  INV_X1 U10438 ( .A(n8044), .ZN(n11665) );
  NAND2_X1 U10439 ( .A1(n11665), .A2(n13056), .ZN(n9137) );
  NAND2_X1 U10440 ( .A1(n9137), .A2(n9135), .ZN(n8046) );
  AOI22_X1 U10441 ( .A1(n12965), .A2(n15195), .B1(n15192), .B2(n13125), .ZN(
        n8047) );
  OAI21_X1 U10442 ( .B1(n8048), .B2(n15198), .A(n8047), .ZN(n13103) );
  NAND2_X1 U10443 ( .A1(n9782), .A2(n12775), .ZN(n15176) );
  NAND2_X1 U10444 ( .A1(n15176), .A2(n15175), .ZN(n15174) );
  NAND2_X1 U10445 ( .A1(n15174), .A2(n12777), .ZN(n10044) );
  NAND2_X1 U10446 ( .A1(n10044), .A2(n12929), .ZN(n10043) );
  NAND2_X1 U10447 ( .A1(n10043), .A2(n12785), .ZN(n10143) );
  NAND2_X1 U10448 ( .A1(n10143), .A2(n12937), .ZN(n10142) );
  NAND2_X1 U10449 ( .A1(n6635), .A2(n10491), .ZN(n12789) );
  NAND2_X1 U10450 ( .A1(n10142), .A2(n12789), .ZN(n10574) );
  NAND2_X1 U10451 ( .A1(n10574), .A2(n12931), .ZN(n8049) );
  NAND2_X1 U10452 ( .A1(n8049), .A2(n12793), .ZN(n10447) );
  NAND2_X1 U10453 ( .A1(n10446), .A2(n12800), .ZN(n10597) );
  INV_X1 U10454 ( .A(n12972), .ZN(n12805) );
  NAND2_X1 U10455 ( .A1(n12805), .A2(n8050), .ZN(n8051) );
  NAND2_X1 U10456 ( .A1(n12970), .A2(n15164), .ZN(n12815) );
  NAND2_X1 U10457 ( .A1(n10995), .A2(n12815), .ZN(n8054) );
  INV_X1 U10458 ( .A(n12970), .ZN(n8053) );
  NAND2_X1 U10459 ( .A1(n8053), .A2(n8052), .ZN(n12816) );
  NAND2_X1 U10460 ( .A1(n8054), .A2(n12816), .ZN(n10878) );
  INV_X1 U10461 ( .A(n10878), .ZN(n8055) );
  XNOR2_X1 U10462 ( .A(n12968), .B(n14769), .ZN(n14772) );
  NAND2_X1 U10463 ( .A1(n12700), .A2(n8057), .ZN(n12827) );
  INV_X1 U10464 ( .A(n12831), .ZN(n8058) );
  AOI21_X2 U10465 ( .B1(n11093), .B2(n12938), .A(n8058), .ZN(n14757) );
  OR2_X1 U10466 ( .A1(n14755), .A2(n13262), .ZN(n12837) );
  AND2_X1 U10467 ( .A1(n14755), .A2(n13262), .ZN(n12839) );
  OR2_X1 U10468 ( .A1(n12736), .A2(n13235), .ZN(n12847) );
  NAND2_X1 U10469 ( .A1(n12736), .A2(n13235), .ZN(n12852) );
  NAND2_X1 U10470 ( .A1(n12847), .A2(n12852), .ZN(n13249) );
  NAND2_X1 U10471 ( .A1(n13236), .A2(n12853), .ZN(n13226) );
  INV_X1 U10472 ( .A(n12858), .ZN(n8059) );
  AOI21_X1 U10473 ( .B1(n13196), .B2(n12869), .A(n8060), .ZN(n13189) );
  NAND2_X1 U10474 ( .A1(n12872), .A2(n13163), .ZN(n12877) );
  NAND2_X1 U10475 ( .A1(n13147), .A2(n13148), .ZN(n13146) );
  XNOR2_X1 U10476 ( .A(n13289), .B(n13151), .ZN(n13140) );
  OR2_X1 U10477 ( .A1(n13289), .A2(n13151), .ZN(n12766) );
  NAND2_X1 U10478 ( .A1(n13107), .A2(n12893), .ZN(n8062) );
  NAND2_X1 U10479 ( .A1(n12564), .A2(n12565), .ZN(n12894) );
  NAND2_X1 U10480 ( .A1(n8062), .A2(n12894), .ZN(n11655) );
  XOR2_X1 U10481 ( .A(n12947), .B(n11655), .Z(n13105) );
  NAND2_X1 U10482 ( .A1(n10042), .A2(n9775), .ZN(n8063) );
  XNOR2_X1 U10483 ( .A(n12962), .B(n8063), .ZN(n8064) );
  AOI21_X1 U10484 ( .B1(n9776), .B2(n10042), .A(n8064), .ZN(n9665) );
  NAND2_X1 U10485 ( .A1(n9776), .A2(n9775), .ZN(n12762) );
  OR3_X1 U10486 ( .A1(n9665), .A2(n13311), .A3(n12762), .ZN(n8066) );
  NOR2_X1 U10487 ( .A1(n12962), .A2(n9775), .ZN(n8065) );
  NAND2_X1 U10488 ( .A1(n9776), .A2(n8065), .ZN(n8110) );
  OR2_X1 U10489 ( .A1(n15200), .A2(n9830), .ZN(n15228) );
  NOR2_X1 U10490 ( .A1(n13105), .A2(n14790), .ZN(n8067) );
  NOR2_X2 U10491 ( .A1(n8068), .A2(P3_IR_REG_22__SCAN_IN), .ZN(n8102) );
  NAND2_X1 U10492 ( .A1(n8102), .A2(n8104), .ZN(n8071) );
  INV_X1 U10493 ( .A(n8071), .ZN(n8070) );
  INV_X1 U10494 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8069) );
  NAND2_X1 U10495 ( .A1(n8070), .A2(n8069), .ZN(n8074) );
  NAND2_X1 U10496 ( .A1(n8071), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8072) );
  XNOR2_X1 U10497 ( .A(n8084), .B(P3_B_REG_SCAN_IN), .ZN(n8077) );
  NAND2_X1 U10498 ( .A1(n8074), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8075) );
  MUX2_X1 U10499 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8075), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8076) );
  NAND2_X1 U10500 ( .A1(n8076), .A2(n6527), .ZN(n10805) );
  NAND2_X1 U10501 ( .A1(n8077), .A2(n10805), .ZN(n8079) );
  NAND2_X1 U10502 ( .A1(n6527), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8078) );
  NAND2_X1 U10503 ( .A1(n8079), .A2(n8086), .ZN(n8087) );
  INV_X1 U10504 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8081) );
  NAND2_X1 U10505 ( .A1(n8899), .A2(n8081), .ZN(n8083) );
  NAND2_X1 U10506 ( .A1(n10805), .A2(n10809), .ZN(n8082) );
  INV_X1 U10507 ( .A(n11777), .ZN(n8085) );
  OAI22_X1 U10508 ( .A1(n8087), .A2(P3_D_REG_0__SCAN_IN), .B1(n8086), .B2(
        n8085), .ZN(n9774) );
  INV_X1 U10509 ( .A(n8089), .ZN(n13388) );
  INV_X1 U10510 ( .A(n13386), .ZN(n8088) );
  NAND2_X1 U10511 ( .A1(n8089), .A2(n8088), .ZN(n8122) );
  INV_X1 U10512 ( .A(n8122), .ZN(n8107) );
  NOR2_X1 U10513 ( .A1(P3_D_REG_10__SCAN_IN), .A2(P3_D_REG_7__SCAN_IN), .ZN(
        n8093) );
  NOR4_X1 U10514 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_2__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n8092) );
  NOR4_X1 U10515 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n8091) );
  NOR4_X1 U10516 ( .A1(P3_D_REG_22__SCAN_IN), .A2(P3_D_REG_25__SCAN_IN), .A3(
        P3_D_REG_20__SCAN_IN), .A4(P3_D_REG_19__SCAN_IN), .ZN(n8090) );
  NAND4_X1 U10517 ( .A1(n8093), .A2(n8092), .A3(n8091), .A4(n8090), .ZN(n8099)
         );
  NOR4_X1 U10518 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n8097) );
  NOR4_X1 U10519 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n8096) );
  NOR4_X1 U10520 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n8095) );
  NOR4_X1 U10521 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n8094) );
  NAND4_X1 U10522 ( .A1(n8097), .A2(n8096), .A3(n8095), .A4(n8094), .ZN(n8098)
         );
  INV_X1 U10523 ( .A(n10805), .ZN(n8101) );
  NOR2_X1 U10524 ( .A1(n11777), .A2(n10809), .ZN(n8100) );
  INV_X1 U10525 ( .A(n8102), .ZN(n8103) );
  INV_X1 U10526 ( .A(n9672), .ZN(n9657) );
  NAND2_X1 U10527 ( .A1(n8120), .A2(n9657), .ZN(n8106) );
  NAND2_X1 U10528 ( .A1(n9776), .A2(n9830), .ZN(n8108) );
  OAI21_X1 U10529 ( .B1(n8117), .B2(n15226), .A(n8108), .ZN(n8109) );
  AOI21_X1 U10530 ( .B1(n8109), .B2(n12762), .A(n12917), .ZN(n8112) );
  NAND2_X1 U10531 ( .A1(n12762), .A2(n12917), .ZN(n9659) );
  NAND2_X1 U10532 ( .A1(n8110), .A2(n12919), .ZN(n9794) );
  NAND2_X1 U10533 ( .A1(n9659), .A2(n9794), .ZN(n9793) );
  NAND2_X1 U10534 ( .A1(n13386), .A2(n9793), .ZN(n8111) );
  OAI21_X1 U10535 ( .B1(n13386), .B2(n8112), .A(n8111), .ZN(n8113) );
  INV_X1 U10536 ( .A(n8114), .ZN(n8115) );
  NAND2_X1 U10537 ( .A1(n10042), .A2(n8117), .ZN(n12954) );
  INV_X1 U10538 ( .A(n12954), .ZN(n8118) );
  AND2_X1 U10539 ( .A1(n8119), .A2(n8118), .ZN(n9663) );
  INV_X1 U10540 ( .A(n9663), .ZN(n9655) );
  INV_X1 U10541 ( .A(n8120), .ZN(n8121) );
  OAI22_X1 U10542 ( .A1(n9671), .A2(n9655), .B1(n9787), .B2(n9665), .ZN(n8123)
         );
  NAND2_X1 U10543 ( .A1(n8123), .A2(n9657), .ZN(n8126) );
  NOR2_X1 U10544 ( .A1(n9672), .A2(n12762), .ZN(n9786) );
  AND2_X1 U10545 ( .A1(n9786), .A2(n12917), .ZN(n9668) );
  INV_X1 U10546 ( .A(n9668), .ZN(n8124) );
  OR2_X1 U10547 ( .A1(n9671), .A2(n8124), .ZN(n8125) );
  INV_X1 U10548 ( .A(n8128), .ZN(n8129) );
  AND3_X2 U10549 ( .A1(n8134), .A2(n8133), .A3(n9406), .ZN(n9544) );
  INV_X1 U10550 ( .A(n8488), .ZN(n8141) );
  NOR2_X1 U10551 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n8146) );
  NAND2_X1 U10552 ( .A1(n8147), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8148) );
  MUX2_X1 U10553 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8148), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8149) );
  NAND2_X1 U10554 ( .A1(n6555), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8150) );
  NOR2_X1 U10555 ( .A1(n14084), .A2(n14089), .ZN(n8151) );
  NAND2_X1 U10556 ( .A1(n11165), .A2(n8151), .ZN(n9093) );
  OR2_X1 U10557 ( .A1(n8153), .A2(n8152), .ZN(n8154) );
  NAND2_X1 U10558 ( .A1(n8155), .A2(n8154), .ZN(n10826) );
  INV_X1 U10559 ( .A(n8578), .ZN(n8156) );
  INV_X1 U10560 ( .A(n8635), .ZN(n8159) );
  NOR2_X1 U10561 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .ZN(n8158) );
  NOR2_X2 U10562 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n9416) );
  NOR2_X2 U10563 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), 
        .ZN(n8161) );
  INV_X1 U10564 ( .A(n8320), .ZN(n8169) );
  NAND2_X1 U10565 ( .A1(n8169), .A2(n8168), .ZN(n8184) );
  INV_X1 U10566 ( .A(n8170), .ZN(n8171) );
  INV_X1 U10567 ( .A(n8180), .ZN(n8172) );
  NOR2_X1 U10568 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .ZN(n8179) );
  NAND2_X1 U10569 ( .A1(n8182), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8183) );
  NAND2_X1 U10570 ( .A1(n8184), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8186) );
  INV_X1 U10571 ( .A(n8348), .ZN(n8187) );
  INV_X1 U10572 ( .A(n9190), .ZN(n9375) );
  INV_X2 U10573 ( .A(n13393), .ZN(n12508) );
  INV_X1 U10574 ( .A(n8188), .ZN(n8190) );
  INV_X1 U10575 ( .A(SI_4_), .ZN(n8189) );
  OAI222_X1 U10576 ( .A1(n9375), .A2(P3_U3151), .B1(n12508), .B2(n8190), .C1(
        n8189), .C2(n9579), .ZN(P3_U3291) );
  INV_X1 U10577 ( .A(n9384), .ZN(n9967) );
  INV_X1 U10578 ( .A(n8191), .ZN(n8193) );
  INV_X1 U10579 ( .A(SI_5_), .ZN(n8192) );
  OAI222_X1 U10580 ( .A1(n9967), .A2(P3_U3151), .B1(n12508), .B2(n8193), .C1(
        n8192), .C2(n9579), .ZN(P3_U3290) );
  OAI222_X1 U10581 ( .A1(P3_U3151), .A2(n15127), .B1(n12508), .B2(n8195), .C1(
        n8194), .C2(n9579), .ZN(P3_U3289) );
  INV_X1 U10582 ( .A(n9478), .ZN(n9179) );
  INV_X1 U10583 ( .A(n8196), .ZN(n8198) );
  INV_X1 U10584 ( .A(SI_3_), .ZN(n8197) );
  OAI222_X1 U10585 ( .A1(n9179), .A2(P3_U3151), .B1(n12508), .B2(n8198), .C1(
        n8197), .C2(n9579), .ZN(P3_U3292) );
  INV_X1 U10586 ( .A(n8199), .ZN(n8201) );
  INV_X1 U10587 ( .A(SI_7_), .ZN(n8200) );
  OAI222_X1 U10588 ( .A1(n10164), .A2(P3_U3151), .B1(n12508), .B2(n8201), .C1(
        n8200), .C2(n9579), .ZN(P3_U3288) );
  INV_X1 U10589 ( .A(n9207), .ZN(n9177) );
  INV_X1 U10590 ( .A(n8202), .ZN(n8203) );
  INV_X1 U10591 ( .A(SI_2_), .ZN(n8219) );
  OAI222_X1 U10592 ( .A1(n9177), .A2(P3_U3151), .B1(n12508), .B2(n8203), .C1(
        n8219), .C2(n9579), .ZN(P3_U3293) );
  NOR2_X1 U10593 ( .A1(n11907), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14070) );
  INV_X2 U10594 ( .A(n14070), .ZN(n14086) );
  INV_X1 U10595 ( .A(n8206), .ZN(n8207) );
  INV_X1 U10596 ( .A(SI_1_), .ZN(n8266) );
  NAND2_X1 U10597 ( .A1(n8232), .A2(n8231), .ZN(n8211) );
  INV_X1 U10598 ( .A(n8211), .ZN(n8209) );
  NAND2_X1 U10599 ( .A1(n8209), .A2(n8230), .ZN(n8218) );
  INV_X1 U10600 ( .A(n8230), .ZN(n8210) );
  NAND2_X1 U10601 ( .A1(n8211), .A2(n8210), .ZN(n8212) );
  NAND2_X1 U10602 ( .A1(n8218), .A2(n8212), .ZN(n8969) );
  NAND2_X1 U10603 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8213) );
  MUX2_X1 U10604 ( .A(n8213), .B(P2_IR_REG_31__SCAN_IN), .S(n13632), .Z(n8215)
         );
  OAI222_X1 U10605 ( .A1(n14086), .A2(n8669), .B1(n14088), .B2(n8969), .C1(
        n8672), .C2(P2_U3088), .ZN(P2_U3326) );
  NAND2_X1 U10606 ( .A1(n8214), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8216) );
  MUX2_X1 U10607 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8216), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n8217) );
  OR2_X1 U10608 ( .A1(n8214), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n8248) );
  NAND2_X1 U10609 ( .A1(n8218), .A2(n8232), .ZN(n8223) );
  INV_X1 U10610 ( .A(n8220), .ZN(n8221) );
  NAND2_X1 U10611 ( .A1(n8233), .A2(n8235), .ZN(n8222) );
  XNOR2_X1 U10612 ( .A(n8223), .B(n8222), .ZN(n8990) );
  INV_X1 U10613 ( .A(n8990), .ZN(n8341) );
  OAI222_X1 U10614 ( .A1(n14992), .A2(P2_U3088), .B1(n14088), .B2(n8341), .C1(
        n8846), .C2(n14086), .ZN(P2_U3325) );
  INV_X1 U10615 ( .A(n8248), .ZN(n8225) );
  INV_X1 U10616 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8224) );
  NAND2_X1 U10617 ( .A1(n8225), .A2(n8224), .ZN(n8250) );
  NAND2_X1 U10618 ( .A1(n8250), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8226) );
  MUX2_X1 U10619 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8226), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8229) );
  INV_X1 U10620 ( .A(n8250), .ZN(n8228) );
  INV_X1 U10621 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8227) );
  NAND2_X1 U10622 ( .A1(n8228), .A2(n8227), .ZN(n8259) );
  INV_X1 U10623 ( .A(n15009), .ZN(n8247) );
  INV_X1 U10624 ( .A(n8232), .ZN(n8234) );
  NAND2_X1 U10625 ( .A1(n8237), .A2(SI_3_), .ZN(n8240) );
  OAI21_X1 U10626 ( .B1(SI_3_), .B2(n8237), .A(n8240), .ZN(n8252) );
  INV_X1 U10627 ( .A(n8252), .ZN(n8238) );
  NAND2_X1 U10628 ( .A1(n8239), .A2(n8238), .ZN(n8254) );
  NAND2_X1 U10629 ( .A1(n8254), .A2(n8240), .ZN(n8242) );
  NAND2_X1 U10630 ( .A1(n8242), .A2(n8241), .ZN(n8257) );
  NAND2_X1 U10631 ( .A1(n8244), .A2(n8243), .ZN(n8245) );
  AND2_X1 U10632 ( .A1(n8257), .A2(n8245), .ZN(n9238) );
  INV_X1 U10633 ( .A(n9238), .ZN(n8295) );
  OAI222_X1 U10634 ( .A1(P2_U3088), .A2(n8247), .B1(n14086), .B2(n8246), .C1(
        n14088), .C2(n8295), .ZN(P2_U3323) );
  NAND2_X1 U10635 ( .A1(n8248), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8249) );
  MUX2_X1 U10636 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8249), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8251) );
  NAND2_X1 U10637 ( .A1(n8253), .A2(n8252), .ZN(n8255) );
  NAND2_X1 U10638 ( .A1(n8255), .A2(n8254), .ZN(n9217) );
  OAI222_X1 U10639 ( .A1(P2_U3088), .A2(n8849), .B1(n14086), .B2(n8850), .C1(
        n14088), .C2(n9217), .ZN(P2_U3324) );
  NAND2_X1 U10640 ( .A1(n8258), .A2(SI_5_), .ZN(n8278) );
  OAI21_X1 U10641 ( .B1(SI_5_), .B2(n8258), .A(n8278), .ZN(n8275) );
  XNOR2_X1 U10642 ( .A(n8277), .B(n8275), .ZN(n9302) );
  INV_X1 U10643 ( .A(n9302), .ZN(n8335) );
  NAND2_X1 U10644 ( .A1(n14070), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8265) );
  NAND2_X1 U10645 ( .A1(n8259), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8260) );
  MUX2_X1 U10646 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8260), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n8264) );
  INV_X1 U10647 ( .A(n8214), .ZN(n8262) );
  INV_X1 U10648 ( .A(n8837), .ZN(n8263) );
  NAND2_X1 U10649 ( .A1(n8935), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15022) );
  OAI211_X1 U10650 ( .C1(n8335), .C2(n14088), .A(n8265), .B(n15022), .ZN(
        P2_U3322) );
  OAI222_X1 U10651 ( .A1(n9173), .A2(P3_U3151), .B1(n12508), .B2(n8267), .C1(
        n8266), .C2(n9579), .ZN(P3_U3294) );
  INV_X1 U10652 ( .A(n8268), .ZN(n8270) );
  INV_X1 U10653 ( .A(SI_9_), .ZN(n8269) );
  OAI222_X1 U10654 ( .A1(n10343), .A2(P3_U3151), .B1(n12508), .B2(n8270), .C1(
        n8269), .C2(n9579), .ZN(P3_U3286) );
  OAI222_X1 U10655 ( .A1(n12508), .A2(n8272), .B1(n9579), .B2(n8271), .C1(
        P3_U3151), .C2(n15149), .ZN(P3_U3287) );
  INV_X1 U10656 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n9159) );
  OAI222_X1 U10657 ( .A1(n12508), .A2(n8273), .B1(P3_U3151), .B2(n9159), .C1(
        n8705), .C2(n9579), .ZN(P3_U3295) );
  OR2_X1 U10658 ( .A1(n8837), .A2(n14068), .ZN(n8274) );
  XNOR2_X1 U10659 ( .A(n8274), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9338) );
  INV_X1 U10660 ( .A(n9338), .ZN(n8286) );
  INV_X1 U10661 ( .A(n8275), .ZN(n8276) );
  NAND2_X1 U10662 ( .A1(n8277), .A2(n8276), .ZN(n8279) );
  NAND2_X1 U10663 ( .A1(n8279), .A2(n8278), .ZN(n8283) );
  MUX2_X1 U10664 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n11907), .Z(n8280) );
  NAND2_X1 U10665 ( .A1(n8280), .A2(SI_6_), .ZN(n8299) );
  OAI21_X1 U10666 ( .B1(SI_6_), .B2(n8280), .A(n8299), .ZN(n8281) );
  INV_X1 U10667 ( .A(n8281), .ZN(n8282) );
  NAND2_X1 U10668 ( .A1(n8283), .A2(n8282), .ZN(n8300) );
  OR2_X1 U10669 ( .A1(n8283), .A2(n8282), .ZN(n8284) );
  AND2_X1 U10670 ( .A1(n8300), .A2(n8284), .ZN(n9616) );
  INV_X1 U10671 ( .A(n9616), .ZN(n8307) );
  OAI222_X1 U10672 ( .A1(P2_U3088), .A2(n8286), .B1(n14086), .B2(n8285), .C1(
        n14088), .C2(n8307), .ZN(P2_U3321) );
  INV_X1 U10673 ( .A(n10346), .ZN(n10508) );
  INV_X1 U10674 ( .A(n8287), .ZN(n8289) );
  INV_X1 U10675 ( .A(SI_10_), .ZN(n8288) );
  OAI222_X1 U10676 ( .A1(n10508), .A2(P3_U3151), .B1(n12508), .B2(n8289), .C1(
        n8288), .C2(n9579), .ZN(P3_U3285) );
  INV_X1 U10677 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8290) );
  NAND2_X1 U10678 ( .A1(n8336), .A2(n8290), .ZN(n8338) );
  OR2_X1 U10679 ( .A1(n8338), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n8310) );
  NAND2_X1 U10680 ( .A1(n8310), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8291) );
  MUX2_X1 U10681 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8291), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n8294) );
  INV_X1 U10682 ( .A(n8310), .ZN(n8293) );
  INV_X1 U10683 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8292) );
  NAND2_X1 U10684 ( .A1(n8293), .A2(n8292), .ZN(n8332) );
  NAND2_X1 U10685 ( .A1(n8294), .A2(n8332), .ZN(n8731) );
  NAND2_X1 U10686 ( .A1(n11907), .A2(P1_U3086), .ZN(n14689) );
  OAI222_X1 U10687 ( .A1(n8731), .A2(P1_U3086), .B1(n14689), .B2(n8296), .C1(
        n14694), .C2(n8295), .ZN(P1_U3351) );
  INV_X1 U10688 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8297) );
  NAND2_X1 U10689 ( .A1(n9422), .A2(n8297), .ZN(n8298) );
  NAND2_X1 U10690 ( .A1(n8298), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8363) );
  XNOR2_X1 U10691 ( .A(n8363), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9926) );
  INV_X1 U10692 ( .A(n9926), .ZN(n8440) );
  NAND2_X1 U10693 ( .A1(n8300), .A2(n8299), .ZN(n8304) );
  MUX2_X1 U10694 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n11907), .Z(n8301) );
  NAND2_X1 U10695 ( .A1(n8301), .A2(SI_7_), .ZN(n8349) );
  OAI21_X1 U10696 ( .B1(SI_7_), .B2(n8301), .A(n8349), .ZN(n8302) );
  INV_X1 U10697 ( .A(n8302), .ZN(n8303) );
  NAND2_X1 U10698 ( .A1(n8304), .A2(n8303), .ZN(n8350) );
  OR2_X1 U10699 ( .A1(n8304), .A2(n8303), .ZN(n8305) );
  OAI222_X1 U10700 ( .A1(n8440), .A2(P1_U3086), .B1(n14689), .B2(n13735), .C1(
        n14694), .C2(n9925), .ZN(P1_U3348) );
  INV_X1 U10701 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14676) );
  OR2_X1 U10702 ( .A1(n9422), .A2(n14676), .ZN(n8306) );
  XNOR2_X1 U10703 ( .A(n8306), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9617) );
  INV_X1 U10704 ( .A(n9617), .ZN(n8414) );
  OAI222_X1 U10705 ( .A1(n8414), .A2(P1_U3086), .B1(n14689), .B2(n8308), .C1(
        n14694), .C2(n8307), .ZN(P1_U3349) );
  NAND2_X1 U10706 ( .A1(n8338), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8309) );
  MUX2_X1 U10707 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8309), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n8311) );
  AND2_X1 U10708 ( .A1(n8311), .A2(n8310), .ZN(n9218) );
  OAI222_X1 U10709 ( .A1(n6865), .A2(P1_U3086), .B1(n14689), .B2(n9219), .C1(
        n14694), .C2(n9217), .ZN(P1_U3352) );
  NAND2_X1 U10710 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8312) );
  MUX2_X1 U10711 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8312), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n8313) );
  NAND2_X1 U10712 ( .A1(n8313), .A2(n7079), .ZN(n14274) );
  INV_X1 U10713 ( .A(n14689), .ZN(n14691) );
  INV_X1 U10714 ( .A(n14691), .ZN(n14684) );
  OAI222_X1 U10715 ( .A1(n14274), .A2(P1_U3086), .B1(n14684), .B2(n8204), .C1(
        n14694), .C2(n8969), .ZN(P1_U3354) );
  INV_X1 U10716 ( .A(n8314), .ZN(n8315) );
  OAI222_X1 U10717 ( .A1(P3_U3151), .A2(n10789), .B1(n12508), .B2(n8315), .C1(
        n8830), .C2(n9579), .ZN(P3_U3284) );
  INV_X1 U10718 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8316) );
  NAND2_X1 U10719 ( .A1(n8837), .A2(n8316), .ZN(n8356) );
  NAND2_X1 U10720 ( .A1(n8356), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8317) );
  XNOR2_X1 U10721 ( .A(n8317), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9432) );
  INV_X1 U10722 ( .A(n9432), .ZN(n8541) );
  INV_X1 U10723 ( .A(n14088), .ZN(n14078) );
  OAI222_X1 U10724 ( .A1(P2_U3088), .A2(n8541), .B1(n14086), .B2(n8318), .C1(
        n14088), .C2(n9925), .ZN(P2_U3320) );
  INV_X1 U10725 ( .A(n8805), .ZN(n8810) );
  INV_X1 U10726 ( .A(n8330), .ZN(n8319) );
  NAND2_X1 U10727 ( .A1(n8319), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12178) );
  NAND2_X1 U10728 ( .A1(n8810), .A2(n12178), .ZN(n8386) );
  NAND2_X1 U10729 ( .A1(n8322), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8324) );
  NAND2_X1 U10730 ( .A1(n8784), .A2(n8710), .ZN(n11927) );
  INV_X1 U10731 ( .A(n11927), .ZN(n9003) );
  XNOR2_X1 U10732 ( .A(n8328), .B(n8327), .ZN(n14683) );
  AOI21_X1 U10733 ( .B1(n9003), .B2(n8330), .A(n11366), .ZN(n8385) );
  INV_X1 U10734 ( .A(n8385), .ZN(n8331) );
  AND2_X1 U10735 ( .A1(n8386), .A2(n8331), .ZN(n14891) );
  NOR2_X1 U10736 ( .A1(n14891), .A2(P1_U4016), .ZN(P1_U3085) );
  NAND2_X1 U10737 ( .A1(n8332), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8333) );
  XNOR2_X1 U10738 ( .A(n8333), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9303) );
  INV_X1 U10739 ( .A(n9303), .ZN(n8401) );
  OAI222_X1 U10740 ( .A1(P1_U3086), .A2(n8401), .B1(n14694), .B2(n8335), .C1(
        n8334), .C2(n14684), .ZN(P1_U3350) );
  NOR2_X1 U10741 ( .A1(n8336), .A2(n14676), .ZN(n8337) );
  MUX2_X1 U10742 ( .A(n14676), .B(n8337), .S(P1_IR_REG_2__SCAN_IN), .Z(n8340)
         );
  INV_X1 U10743 ( .A(n8338), .ZN(n8339) );
  NOR2_X1 U10744 ( .A1(n8340), .A2(n8339), .ZN(n8991) );
  OAI222_X1 U10745 ( .A1(P1_U3086), .A2(n7065), .B1(n14694), .B2(n8341), .C1(
        n13734), .C2(n14684), .ZN(P1_U3353) );
  INV_X1 U10746 ( .A(P1_B_REG_SCAN_IN), .ZN(n11463) );
  NOR2_X1 U10747 ( .A1(n14692), .A2(n11463), .ZN(n8342) );
  NAND2_X1 U10748 ( .A1(n11164), .A2(n8342), .ZN(n8343) );
  INV_X1 U10749 ( .A(n8780), .ZN(n8345) );
  NAND2_X1 U10750 ( .A1(n8345), .A2(n8805), .ZN(n14917) );
  INV_X1 U10751 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n8779) );
  INV_X1 U10752 ( .A(n8347), .ZN(n14690) );
  AND2_X1 U10753 ( .A1(n8348), .A2(n14690), .ZN(n8346) );
  AOI22_X1 U10754 ( .A1(n14917), .A2(n8779), .B1(n8346), .B2(n11164), .ZN(
        P1_U3445) );
  INV_X1 U10755 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n8776) );
  NOR2_X1 U10756 ( .A1(n14692), .A2(n8347), .ZN(n8775) );
  AOI22_X1 U10757 ( .A1(n14917), .A2(n8776), .B1(n8348), .B2(n8775), .ZN(
        P1_U3446) );
  MUX2_X1 U10758 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n11907), .Z(n8351) );
  NAND2_X1 U10759 ( .A1(n8351), .A2(SI_8_), .ZN(n8371) );
  OAI21_X1 U10760 ( .B1(SI_8_), .B2(n8351), .A(n8371), .ZN(n8352) );
  INV_X1 U10761 ( .A(n8352), .ZN(n8353) );
  NAND2_X1 U10762 ( .A1(n8359), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8357) );
  MUX2_X1 U10763 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8357), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n8358) );
  INV_X1 U10764 ( .A(n8358), .ZN(n8360) );
  NOR2_X1 U10765 ( .A1(n8359), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8378) );
  NOR2_X1 U10766 ( .A1(n8360), .A2(n8378), .ZN(n9483) );
  NAND2_X1 U10767 ( .A1(n9483), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15033) );
  NAND2_X1 U10768 ( .A1(n14070), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8361) );
  OAI211_X1 U10769 ( .C1(n10098), .C2(n14088), .A(n15033), .B(n8361), .ZN(
        P2_U3319) );
  OAI222_X1 U10770 ( .A1(n9579), .A2(n9029), .B1(n12508), .B2(n8362), .C1(
        n12985), .C2(P3_U3151), .ZN(P3_U3283) );
  NAND2_X1 U10771 ( .A1(n8363), .A2(n9417), .ZN(n8364) );
  NAND2_X1 U10772 ( .A1(n8364), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8637) );
  XNOR2_X1 U10773 ( .A(n8637), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10099) );
  INV_X1 U10774 ( .A(n10099), .ZN(n8448) );
  OAI222_X1 U10775 ( .A1(n8448), .A2(P1_U3086), .B1(n14689), .B2(n8365), .C1(
        n14694), .C2(n10098), .ZN(P1_U3347) );
  NAND2_X1 U10776 ( .A1(n8637), .A2(n8366), .ZN(n8367) );
  NAND2_X1 U10777 ( .A1(n8367), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8369) );
  NAND2_X1 U10778 ( .A1(n8369), .A2(n8368), .ZN(n8470) );
  OR2_X1 U10779 ( .A1(n8369), .A2(n8368), .ZN(n8370) );
  INV_X1 U10780 ( .A(n10380), .ZN(n8456) );
  MUX2_X1 U10781 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n11907), .Z(n8373) );
  NAND2_X1 U10782 ( .A1(n8373), .A2(SI_9_), .ZN(n8462) );
  OAI21_X1 U10783 ( .B1(SI_9_), .B2(n8373), .A(n8462), .ZN(n8374) );
  INV_X1 U10784 ( .A(n8374), .ZN(n8375) );
  OAI222_X1 U10785 ( .A1(n8456), .A2(P1_U3086), .B1(n14689), .B2(n8377), .C1(
        n14694), .C2(n10379), .ZN(P1_U3346) );
  INV_X1 U10786 ( .A(n8378), .ZN(n8380) );
  NAND2_X1 U10787 ( .A1(n8380), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8379) );
  MUX2_X1 U10788 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8379), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n8381) );
  INV_X1 U10789 ( .A(n9705), .ZN(n8524) );
  OAI222_X1 U10790 ( .A1(P2_U3088), .A2(n8524), .B1(n14086), .B2(n8382), .C1(
        n14088), .C2(n10379), .ZN(P2_U3318) );
  OAI222_X1 U10791 ( .A1(n11127), .A2(P3_U3151), .B1(n12508), .B2(n8383), .C1(
        n9033), .C2(n9579), .ZN(P3_U3282) );
  NAND2_X1 U10792 ( .A1(n8386), .A2(n8385), .ZN(n14894) );
  INV_X1 U10793 ( .A(n14683), .ZN(n9002) );
  INV_X1 U10794 ( .A(n6663), .ZN(n12174) );
  OR2_X1 U10795 ( .A1(n14894), .A2(n12174), .ZN(n14323) );
  INV_X1 U10796 ( .A(n14323), .ZN(n14901) );
  INV_X1 U10797 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9254) );
  XNOR2_X1 U10798 ( .A(n9303), .B(n9254), .ZN(n8388) );
  INV_X1 U10799 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n8997) );
  INV_X1 U10800 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n8986) );
  MUX2_X1 U10801 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n8986), .S(n8991), .Z(n8738)
         );
  INV_X1 U10802 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n8788) );
  MUX2_X1 U10803 ( .A(n8788), .B(P1_REG1_REG_1__SCAN_IN), .S(n14274), .Z(
        n14270) );
  AND2_X1 U10804 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14269) );
  NAND2_X1 U10805 ( .A1(n14270), .A2(n14269), .ZN(n14268) );
  OAI21_X1 U10806 ( .B1(n14274), .B2(n8788), .A(n14268), .ZN(n8737) );
  NAND2_X1 U10807 ( .A1(n8738), .A2(n8737), .ZN(n8736) );
  OAI21_X1 U10808 ( .B1(n7065), .B2(n8986), .A(n8736), .ZN(n14283) );
  MUX2_X1 U10809 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n8997), .S(n9218), .Z(n14284) );
  NAND2_X1 U10810 ( .A1(n14283), .A2(n14284), .ZN(n14282) );
  OAI21_X1 U10811 ( .B1(n8997), .B2(n6865), .A(n14282), .ZN(n8719) );
  INV_X1 U10812 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9468) );
  MUX2_X1 U10813 ( .A(n9468), .B(P1_REG1_REG_4__SCAN_IN), .S(n8731), .Z(n8720)
         );
  INV_X1 U10814 ( .A(n8731), .ZN(n9239) );
  AOI22_X1 U10815 ( .A1(n8719), .A2(n8720), .B1(n9239), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n8387) );
  NAND2_X1 U10816 ( .A1(n8387), .A2(n8388), .ZN(n8402) );
  OAI21_X1 U10817 ( .B1(n8388), .B2(n8387), .A(n8402), .ZN(n8397) );
  NAND2_X1 U10818 ( .A1(n9002), .A2(n12174), .ZN(n8389) );
  INV_X1 U10819 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n8983) );
  MUX2_X1 U10820 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n8983), .S(n8991), .Z(n8735)
         );
  INV_X1 U10821 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n8390) );
  MUX2_X1 U10822 ( .A(n8390), .B(P1_REG2_REG_1__SCAN_IN), .S(n14274), .Z(
        n14272) );
  AND2_X1 U10823 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14273) );
  NAND2_X1 U10824 ( .A1(n14272), .A2(n14273), .ZN(n14271) );
  OAI21_X1 U10825 ( .B1(n8390), .B2(n14274), .A(n14271), .ZN(n8734) );
  AND2_X1 U10826 ( .A1(n8735), .A2(n8734), .ZN(n14287) );
  NOR2_X1 U10827 ( .A1(n7065), .A2(n8983), .ZN(n14286) );
  INV_X1 U10828 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9508) );
  MUX2_X1 U10829 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9508), .S(n9218), .Z(n14285) );
  OAI21_X1 U10830 ( .B1(n14287), .B2(n14286), .A(n14285), .ZN(n14289) );
  NAND2_X1 U10831 ( .A1(n9218), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8726) );
  INV_X1 U10832 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n8391) );
  MUX2_X1 U10833 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n8391), .S(n8731), .Z(n8725)
         );
  AOI21_X1 U10834 ( .B1(n14289), .B2(n8726), .A(n8725), .ZN(n8724) );
  NOR2_X1 U10835 ( .A1(n8731), .A2(n8391), .ZN(n8393) );
  INV_X1 U10836 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9688) );
  MUX2_X1 U10837 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9688), .S(n9303), .Z(n8392)
         );
  OAI21_X1 U10838 ( .B1(n8724), .B2(n8393), .A(n8392), .ZN(n8407) );
  INV_X1 U10839 ( .A(n8407), .ZN(n8395) );
  NOR3_X1 U10840 ( .A1(n8724), .A2(n8393), .A3(n8392), .ZN(n8394) );
  NOR3_X1 U10841 ( .A1(n14906), .A2(n8395), .A3(n8394), .ZN(n8396) );
  AOI21_X1 U10842 ( .B1(n14901), .B2(n8397), .A(n8396), .ZN(n8400) );
  NAND2_X1 U10843 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9319) );
  INV_X1 U10844 ( .A(n9319), .ZN(n8398) );
  AOI21_X1 U10845 ( .B1(n14891), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n8398), .ZN(
        n8399) );
  OAI211_X1 U10846 ( .C1(n8401), .C2(n14320), .A(n8400), .B(n8399), .ZN(
        P1_U3248) );
  INV_X1 U10847 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9314) );
  MUX2_X1 U10848 ( .A(n9314), .B(P1_REG1_REG_6__SCAN_IN), .S(n9617), .Z(n8404)
         );
  OAI21_X1 U10849 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n9303), .A(n8402), .ZN(
        n8403) );
  NOR2_X1 U10850 ( .A1(n8403), .A2(n8404), .ZN(n8419) );
  AOI211_X1 U10851 ( .C1(n8404), .C2(n8403), .A(n8419), .B(n14323), .ZN(n8410)
         );
  NAND2_X1 U10852 ( .A1(n9303), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8406) );
  INV_X1 U10853 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n8413) );
  MUX2_X1 U10854 ( .A(n8413), .B(P1_REG2_REG_6__SCAN_IN), .S(n9617), .Z(n8405)
         );
  AOI21_X1 U10855 ( .B1(n8407), .B2(n8406), .A(n8405), .ZN(n8436) );
  AND3_X1 U10856 ( .A1(n8407), .A2(n8406), .A3(n8405), .ZN(n8408) );
  NOR3_X1 U10857 ( .A1(n14906), .A2(n8436), .A3(n8408), .ZN(n8409) );
  NOR2_X1 U10858 ( .A1(n8410), .A2(n8409), .ZN(n8412) );
  AND2_X1 U10859 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9637) );
  AOI21_X1 U10860 ( .B1(n14891), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n9637), .ZN(
        n8411) );
  OAI211_X1 U10861 ( .C1(n8414), .C2(n14320), .A(n8412), .B(n8411), .ZN(
        P1_U3249) );
  NOR2_X1 U10862 ( .A1(n8414), .A2(n8413), .ZN(n8431) );
  INV_X1 U10863 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9949) );
  MUX2_X1 U10864 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9949), .S(n9926), .Z(n8415)
         );
  OAI21_X1 U10865 ( .B1(n8436), .B2(n8431), .A(n8415), .ZN(n8434) );
  NAND2_X1 U10866 ( .A1(n9926), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8417) );
  INV_X1 U10867 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n8447) );
  MUX2_X1 U10868 ( .A(n8447), .B(P1_REG2_REG_8__SCAN_IN), .S(n10099), .Z(n8416) );
  AOI21_X1 U10869 ( .B1(n8434), .B2(n8417), .A(n8416), .ZN(n8451) );
  NAND3_X1 U10870 ( .A1(n8434), .A2(n8417), .A3(n8416), .ZN(n8418) );
  NAND2_X1 U10871 ( .A1(n14318), .A2(n8418), .ZN(n8427) );
  AOI21_X1 U10872 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n9617), .A(n8419), .ZN(
        n8430) );
  INV_X1 U10873 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9631) );
  MUX2_X1 U10874 ( .A(n9631), .B(P1_REG1_REG_7__SCAN_IN), .S(n9926), .Z(n8429)
         );
  NOR2_X1 U10875 ( .A1(n8430), .A2(n8429), .ZN(n8428) );
  AOI21_X1 U10876 ( .B1(n9926), .B2(P1_REG1_REG_7__SCAN_IN), .A(n8428), .ZN(
        n8421) );
  INV_X1 U10877 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9933) );
  MUX2_X1 U10878 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9933), .S(n10099), .Z(n8420) );
  NAND2_X1 U10879 ( .A1(n8421), .A2(n8420), .ZN(n8444) );
  OAI21_X1 U10880 ( .B1(n8421), .B2(n8420), .A(n8444), .ZN(n8422) );
  NAND2_X1 U10881 ( .A1(n8422), .A2(n14901), .ZN(n8426) );
  INV_X1 U10882 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n13634) );
  NOR2_X1 U10883 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13634), .ZN(n8424) );
  NOR2_X1 U10884 ( .A1(n14320), .A2(n8448), .ZN(n8423) );
  AOI211_X1 U10885 ( .C1(n14891), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n8424), .B(
        n8423), .ZN(n8425) );
  OAI211_X1 U10886 ( .C1(n8451), .C2(n8427), .A(n8426), .B(n8425), .ZN(
        P1_U3251) );
  AOI211_X1 U10887 ( .C1(n8430), .C2(n8429), .A(n14323), .B(n8428), .ZN(n8442)
         );
  INV_X1 U10888 ( .A(n8431), .ZN(n8433) );
  MUX2_X1 U10889 ( .A(n9949), .B(P1_REG2_REG_7__SCAN_IN), .S(n9926), .Z(n8432)
         );
  NAND2_X1 U10890 ( .A1(n8433), .A2(n8432), .ZN(n8435) );
  OAI211_X1 U10891 ( .C1(n8436), .C2(n8435), .A(n14318), .B(n8434), .ZN(n8439)
         );
  AND2_X1 U10892 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8437) );
  AOI21_X1 U10893 ( .B1(n14891), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n8437), .ZN(
        n8438) );
  OAI211_X1 U10894 ( .C1(n14320), .C2(n8440), .A(n8439), .B(n8438), .ZN(n8441)
         );
  OR2_X1 U10895 ( .A1(n8442), .A2(n8441), .ZN(P1_U3250) );
  INV_X1 U10896 ( .A(n11122), .ZN(n11134) );
  OAI222_X1 U10897 ( .A1(n9579), .A2(n9413), .B1(n12508), .B2(n8443), .C1(
        n11134), .C2(P3_U3151), .ZN(P3_U3281) );
  INV_X1 U10898 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10119) );
  MUX2_X1 U10899 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10119), .S(n10380), .Z(
        n8446) );
  OAI21_X1 U10900 ( .B1(n10099), .B2(P1_REG1_REG_8__SCAN_IN), .A(n8444), .ZN(
        n8445) );
  NAND2_X1 U10901 ( .A1(n8445), .A2(n8446), .ZN(n8745) );
  OAI21_X1 U10902 ( .B1(n8446), .B2(n8445), .A(n8745), .ZN(n8459) );
  NOR2_X1 U10903 ( .A1(n8448), .A2(n8447), .ZN(n8450) );
  INV_X1 U10904 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10398) );
  MUX2_X1 U10905 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10398), .S(n10380), .Z(
        n8449) );
  OAI21_X1 U10906 ( .B1(n8451), .B2(n8450), .A(n8449), .ZN(n8751) );
  INV_X1 U10907 ( .A(n8751), .ZN(n8453) );
  NOR3_X1 U10908 ( .A1(n8451), .A2(n8450), .A3(n8449), .ZN(n8452) );
  NOR3_X1 U10909 ( .A1(n8453), .A2(n8452), .A3(n14906), .ZN(n8458) );
  NAND2_X1 U10910 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n14880) );
  INV_X1 U10911 ( .A(n14880), .ZN(n8454) );
  AOI21_X1 U10912 ( .B1(n14891), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n8454), .ZN(
        n8455) );
  OAI21_X1 U10913 ( .B1(n14320), .B2(n8456), .A(n8455), .ZN(n8457) );
  AOI211_X1 U10914 ( .C1(n8459), .C2(n14901), .A(n8458), .B(n8457), .ZN(n8460)
         );
  INV_X1 U10915 ( .A(n8460), .ZN(P1_U3252) );
  NAND2_X1 U10916 ( .A1(n8629), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8461) );
  XNOR2_X1 U10917 ( .A(n8461), .B(P2_IR_REG_10__SCAN_IN), .ZN(n9841) );
  INV_X1 U10918 ( .A(n9841), .ZN(n8665) );
  MUX2_X1 U10919 ( .A(n8472), .B(n8469), .S(n11907), .Z(n8466) );
  NAND2_X1 U10920 ( .A1(n8467), .A2(n8466), .ZN(n8468) );
  OAI222_X1 U10921 ( .A1(P2_U3088), .A2(n8665), .B1(n14086), .B2(n8469), .C1(
        n14088), .C2(n10527), .ZN(P2_U3317) );
  NAND2_X1 U10922 ( .A1(n8470), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8471) );
  XNOR2_X1 U10923 ( .A(n8471), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10528) );
  INV_X1 U10924 ( .A(n10528), .ZN(n8755) );
  OAI222_X1 U10925 ( .A1(n8755), .A2(P1_U3086), .B1(n14684), .B2(n8472), .C1(
        n14694), .C2(n10527), .ZN(P1_U3345) );
  INV_X1 U10926 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n8473) );
  MUX2_X1 U10927 ( .A(n8473), .B(P2_REG1_REG_3__SCAN_IN), .S(n8849), .Z(n8623)
         );
  INV_X1 U10928 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n8687) );
  MUX2_X1 U10929 ( .A(n8687), .B(P2_REG1_REG_1__SCAN_IN), .S(n8672), .Z(n8643)
         );
  AND2_X1 U10930 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n8642) );
  NAND2_X1 U10931 ( .A1(n8643), .A2(n8642), .ZN(n8641) );
  INV_X1 U10932 ( .A(n8672), .ZN(n8653) );
  NAND2_X1 U10933 ( .A1(n8653), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8474) );
  NAND2_X1 U10934 ( .A1(n8641), .A2(n8474), .ZN(n14989) );
  INV_X1 U10935 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n8475) );
  MUX2_X1 U10936 ( .A(n8475), .B(P2_REG1_REG_2__SCAN_IN), .S(n14992), .Z(
        n14990) );
  INV_X1 U10937 ( .A(n14992), .ZN(n8506) );
  NAND2_X1 U10938 ( .A1(n8506), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8476) );
  NAND2_X1 U10939 ( .A1(n14988), .A2(n8476), .ZN(n8622) );
  NAND2_X1 U10940 ( .A1(n8623), .A2(n8622), .ZN(n8621) );
  INV_X1 U10941 ( .A(n8849), .ZN(n8477) );
  NAND2_X1 U10942 ( .A1(n8477), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8478) );
  INV_X1 U10943 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n15107) );
  MUX2_X1 U10944 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n15107), .S(n15009), .Z(
        n15005) );
  NAND2_X1 U10945 ( .A1(n15009), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8479) );
  NAND2_X1 U10946 ( .A1(n15002), .A2(n8479), .ZN(n15017) );
  INV_X1 U10947 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n8480) );
  MUX2_X1 U10948 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n8480), .S(n8935), .Z(n15018) );
  NAND2_X1 U10949 ( .A1(n8935), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8481) );
  NAND2_X1 U10950 ( .A1(n15016), .A2(n8481), .ZN(n8556) );
  INV_X1 U10951 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n15110) );
  MUX2_X1 U10952 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n15110), .S(n9338), .Z(n8557) );
  NAND2_X1 U10953 ( .A1(n8556), .A2(n8557), .ZN(n8555) );
  NAND2_X1 U10954 ( .A1(n9338), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8482) );
  NAND2_X1 U10955 ( .A1(n8555), .A2(n8482), .ZN(n8537) );
  INV_X1 U10956 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n8483) );
  MUX2_X1 U10957 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n8483), .S(n9432), .Z(n8538)
         );
  INV_X1 U10958 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n8484) );
  MUX2_X1 U10959 ( .A(n8484), .B(P2_REG1_REG_8__SCAN_IN), .S(n9483), .Z(n15030) );
  NOR2_X1 U10960 ( .A1(n15031), .A2(n15030), .ZN(n15029) );
  INV_X1 U10961 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8485) );
  MUX2_X1 U10962 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n8485), .S(n9705), .Z(n8486)
         );
  NAND2_X1 U10963 ( .A1(n8487), .A2(n8486), .ZN(n8656) );
  OAI21_X1 U10964 ( .B1(n8487), .B2(n8486), .A(n8656), .ZN(n8504) );
  INV_X1 U10965 ( .A(n10826), .ZN(n9091) );
  OR2_X1 U10966 ( .A1(n9093), .A2(n9091), .ZN(n8499) );
  NAND2_X1 U10967 ( .A1(n9117), .A2(n10826), .ZN(n8497) );
  XNOR2_X1 U10968 ( .A(n8494), .B(n8496), .ZN(n8500) );
  NAND2_X1 U10969 ( .A1(n8497), .A2(n8931), .ZN(n8498) );
  AND2_X1 U10970 ( .A1(n8499), .A2(n8498), .ZN(n8522) );
  INV_X1 U10971 ( .A(n8606), .ZN(n8675) );
  NAND2_X1 U10972 ( .A1(n8675), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14079) );
  INV_X1 U10973 ( .A(n14079), .ZN(n8502) );
  AND2_X1 U10974 ( .A1(n8502), .A2(n8501), .ZN(n8503) );
  NAND2_X1 U10975 ( .A1(n8504), .A2(n15003), .ZN(n8528) );
  INV_X1 U10976 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8516) );
  INV_X1 U10977 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n13909) );
  MUX2_X1 U10978 ( .A(n13909), .B(P2_REG2_REG_3__SCAN_IN), .S(n8849), .Z(n8507) );
  INV_X1 U10979 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n13928) );
  MUX2_X1 U10980 ( .A(n13928), .B(P2_REG2_REG_1__SCAN_IN), .S(n8672), .Z(n8645) );
  AND2_X1 U10981 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n8646) );
  NAND2_X1 U10982 ( .A1(n8645), .A2(n8646), .ZN(n8644) );
  NAND2_X1 U10983 ( .A1(n8653), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8505) );
  NAND2_X1 U10984 ( .A1(n8644), .A2(n8505), .ZN(n14997) );
  INV_X1 U10985 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n13917) );
  MUX2_X1 U10986 ( .A(n13917), .B(P2_REG2_REG_2__SCAN_IN), .S(n14992), .Z(
        n14996) );
  NAND2_X1 U10987 ( .A1(n14997), .A2(n14996), .ZN(n14995) );
  NAND2_X1 U10988 ( .A1(n8506), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8615) );
  OR2_X1 U10989 ( .A1(n8849), .A2(n13909), .ZN(n8508) );
  NAND2_X1 U10990 ( .A1(n8618), .A2(n8508), .ZN(n15012) );
  INV_X1 U10991 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10305) );
  MUX2_X1 U10992 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10305), .S(n15009), .Z(
        n15011) );
  NAND2_X1 U10993 ( .A1(n15012), .A2(n15011), .ZN(n15010) );
  NAND2_X1 U10994 ( .A1(n15009), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8509) );
  NAND2_X1 U10995 ( .A1(n15010), .A2(n8509), .ZN(n15026) );
  INV_X1 U10996 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10031) );
  MUX2_X1 U10997 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10031), .S(n8935), .Z(
        n15025) );
  NAND2_X1 U10998 ( .A1(n8935), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8550) );
  NAND2_X1 U10999 ( .A1(n15024), .A2(n8550), .ZN(n8511) );
  INV_X1 U11000 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10317) );
  MUX2_X1 U11001 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10317), .S(n9338), .Z(n8510) );
  NAND2_X1 U11002 ( .A1(n8511), .A2(n8510), .ZN(n8552) );
  NAND2_X1 U11003 ( .A1(n9338), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8530) );
  NAND2_X1 U11004 ( .A1(n8552), .A2(n8530), .ZN(n8514) );
  INV_X1 U11005 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n8512) );
  MUX2_X1 U11006 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n8512), .S(n9432), .Z(n8513)
         );
  NAND2_X1 U11007 ( .A1(n8514), .A2(n8513), .ZN(n8532) );
  NAND2_X1 U11008 ( .A1(n9432), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8515) );
  NAND2_X1 U11009 ( .A1(n8532), .A2(n8515), .ZN(n15041) );
  MUX2_X1 U11010 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n8516), .S(n9483), .Z(n15040) );
  AND2_X1 U11011 ( .A1(n15041), .A2(n15040), .ZN(n15037) );
  INV_X1 U11012 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8517) );
  MUX2_X1 U11013 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n8517), .S(n9705), .Z(n8518)
         );
  NAND2_X1 U11014 ( .A1(n8519), .A2(n8518), .ZN(n8659) );
  OAI21_X1 U11015 ( .B1(n8519), .B2(n8518), .A(n8659), .ZN(n8526) );
  NOR2_X1 U11016 ( .A1(n8501), .A2(n14079), .ZN(n8520) );
  NAND2_X1 U11017 ( .A1(n8521), .A2(n8606), .ZN(n15034) );
  OR2_X1 U11018 ( .A1(n15034), .A2(P2_U3088), .ZN(n14993) );
  AND2_X1 U11019 ( .A1(n8522), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14987) );
  NAND2_X1 U11020 ( .A1(n14987), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U11021 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n9717) );
  OAI211_X1 U11022 ( .C1(n14993), .C2(n8524), .A(n8523), .B(n9717), .ZN(n8525)
         );
  AOI21_X1 U11023 ( .B1(n8526), .B2(n15039), .A(n8525), .ZN(n8527) );
  NAND2_X1 U11024 ( .A1(n8528), .A2(n8527), .ZN(P2_U3223) );
  INV_X1 U11025 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n13710) );
  NOR2_X1 U11026 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13710), .ZN(n8534) );
  MUX2_X1 U11027 ( .A(n8512), .B(P2_REG2_REG_7__SCAN_IN), .S(n9432), .Z(n8529)
         );
  NAND3_X1 U11028 ( .A1(n8552), .A2(n8530), .A3(n8529), .ZN(n8531) );
  AND3_X1 U11029 ( .A1(n15039), .A2(n8532), .A3(n8531), .ZN(n8533) );
  AOI211_X1 U11030 ( .C1(n14987), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n8534), .B(
        n8533), .ZN(n8540) );
  INV_X1 U11031 ( .A(n8535), .ZN(n8536) );
  OAI211_X1 U11032 ( .C1(n8538), .C2(n8537), .A(n15003), .B(n8536), .ZN(n8539)
         );
  OAI211_X1 U11033 ( .C1(n14993), .C2(n8541), .A(n8540), .B(n8539), .ZN(
        P2_U3221) );
  INV_X1 U11034 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n8614) );
  INV_X1 U11035 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n8542) );
  NAND2_X1 U11036 ( .A1(n15039), .A2(n8542), .ZN(n8543) );
  OAI211_X1 U11037 ( .C1(n15046), .C2(P2_REG1_REG_0__SCAN_IN), .A(n8543), .B(
        n14993), .ZN(n8544) );
  INV_X1 U11038 ( .A(n8544), .ZN(n8546) );
  AOI22_X1 U11039 ( .A1(n15003), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n15039), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n8545) );
  INV_X1 U11040 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8600) );
  MUX2_X1 U11041 ( .A(n8546), .B(n8545), .S(n8600), .Z(n8548) );
  AOI22_X1 U11042 ( .A1(n14987), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n8547) );
  NAND2_X1 U11043 ( .A1(n8548), .A2(n8547), .ZN(P2_U3214) );
  INV_X1 U11044 ( .A(n14993), .ZN(n15052) );
  NAND2_X1 U11045 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n9358) );
  INV_X1 U11046 ( .A(n9358), .ZN(n8554) );
  MUX2_X1 U11047 ( .A(n10317), .B(P2_REG2_REG_6__SCAN_IN), .S(n9338), .Z(n8549) );
  NAND3_X1 U11048 ( .A1(n15024), .A2(n8550), .A3(n8549), .ZN(n8551) );
  AND3_X1 U11049 ( .A1(n15039), .A2(n8552), .A3(n8551), .ZN(n8553) );
  AOI211_X1 U11050 ( .C1(n15052), .C2(n9338), .A(n8554), .B(n8553), .ZN(n8559)
         );
  OAI211_X1 U11051 ( .C1(n8557), .C2(n8556), .A(n15003), .B(n8555), .ZN(n8558)
         );
  OAI211_X1 U11052 ( .C1(n7493), .C2(n15061), .A(n8559), .B(n8558), .ZN(
        P2_U3220) );
  INV_X1 U11053 ( .A(n11272), .ZN(n13010) );
  OAI222_X1 U11054 ( .A1(n9579), .A2(n9538), .B1(n12508), .B2(n8560), .C1(
        n13010), .C2(P3_U3151), .ZN(P3_U3280) );
  NOR4_X1 U11055 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n8564) );
  NOR4_X1 U11056 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n8563) );
  NOR4_X1 U11057 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8562) );
  NOR4_X1 U11058 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8561) );
  AND4_X1 U11059 ( .A1(n8564), .A2(n8563), .A3(n8562), .A4(n8561), .ZN(n8572)
         );
  NOR2_X1 U11060 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .ZN(
        n13724) );
  NOR4_X1 U11061 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n8567) );
  NOR4_X1 U11062 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n8566) );
  NOR4_X1 U11063 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n8565) );
  AND4_X1 U11064 ( .A1(n13724), .A2(n8567), .A3(n8566), .A4(n8565), .ZN(n8571)
         );
  XOR2_X1 U11065 ( .A(P2_B_REG_SCAN_IN), .B(n11165), .Z(n8568) );
  INV_X1 U11066 ( .A(n15076), .ZN(n8570) );
  NOR2_X1 U11067 ( .A1(n8573), .A2(n14068), .ZN(n8574) );
  NAND2_X1 U11068 ( .A1(n8575), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8577) );
  NAND2_X1 U11069 ( .A1(n6629), .A2(n13574), .ZN(n12443) );
  AND2_X1 U11070 ( .A1(n12443), .A2(n12441), .ZN(n12404) );
  AND2_X1 U11071 ( .A1(n12404), .A2(n12498), .ZN(n9092) );
  INV_X1 U11072 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15086) );
  NAND2_X1 U11073 ( .A1(n15076), .A2(n15086), .ZN(n8580) );
  NAND2_X1 U11074 ( .A1(n14084), .A2(n14089), .ZN(n8579) );
  NAND2_X1 U11075 ( .A1(n8580), .A2(n8579), .ZN(n9087) );
  NAND3_X1 U11076 ( .A1(n15087), .A2(n9087), .A3(n9099), .ZN(n8581) );
  INV_X1 U11077 ( .A(n14084), .ZN(n8582) );
  OR2_X1 U11078 ( .A1(n11165), .A2(n8582), .ZN(n8584) );
  INV_X1 U11079 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15083) );
  NAND2_X1 U11080 ( .A1(n15076), .A2(n15083), .ZN(n8583) );
  INV_X1 U11081 ( .A(n15084), .ZN(n9125) );
  NAND2_X1 U11082 ( .A1(n12390), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U11083 ( .A1(n8853), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8596) );
  NAND2_X1 U11084 ( .A1(n11528), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8595) );
  NAND2_X1 U11085 ( .A1(n6446), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8594) );
  INV_X1 U11086 ( .A(n12180), .ZN(n12183) );
  NAND2_X1 U11087 ( .A1(n11907), .A2(SI_0_), .ZN(n8599) );
  XNOR2_X1 U11088 ( .A(n8599), .B(n8598), .ZN(n14090) );
  NAND2_X1 U11089 ( .A1(n12183), .A2(n9834), .ZN(n8681) );
  NAND2_X1 U11090 ( .A1(n12185), .A2(n13563), .ZN(n8601) );
  AND2_X1 U11091 ( .A1(n8681), .A2(n8601), .ZN(n12450) );
  NAND2_X1 U11092 ( .A1(n12498), .A2(n13603), .ZN(n8604) );
  INV_X1 U11093 ( .A(n6629), .ZN(n12449) );
  NAND2_X1 U11094 ( .A1(n12449), .A2(n12441), .ZN(n8603) );
  AOI21_X1 U11095 ( .B1(n13875), .B2(n6597), .A(n12450), .ZN(n8612) );
  NAND2_X1 U11096 ( .A1(n9117), .A2(n8606), .ZN(n11617) );
  INV_X2 U11097 ( .A(n11617), .ZN(n13517) );
  NAND2_X1 U11098 ( .A1(n11528), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8610) );
  NAND2_X1 U11099 ( .A1(n6446), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U11100 ( .A1(n8853), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8607) );
  NAND2_X1 U11101 ( .A1(n13517), .A2(n13561), .ZN(n9840) );
  INV_X1 U11102 ( .A(n9840), .ZN(n8611) );
  NOR2_X1 U11103 ( .A1(n8612), .A2(n8611), .ZN(n9129) );
  NAND3_X1 U11104 ( .A1(n9834), .A2(n12179), .A3(n6667), .ZN(n9130) );
  OAI211_X1 U11105 ( .C1(n12450), .C2(n15101), .A(n9129), .B(n9130), .ZN(n8799) );
  NAND2_X1 U11106 ( .A1(n15112), .A2(n8799), .ZN(n8613) );
  OAI21_X1 U11107 ( .B1(n15112), .B2(n8614), .A(n8613), .ZN(P2_U3499) );
  INV_X1 U11108 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n8620) );
  MUX2_X1 U11109 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n13909), .S(n8849), .Z(n8616) );
  NAND3_X1 U11110 ( .A1(n8616), .A2(n14995), .A3(n8615), .ZN(n8617) );
  NAND3_X1 U11111 ( .A1(n15039), .A2(n8618), .A3(n8617), .ZN(n8619) );
  OAI21_X1 U11112 ( .B1(n15061), .B2(n8620), .A(n8619), .ZN(n8627) );
  INV_X1 U11113 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9097) );
  NOR2_X1 U11114 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9097), .ZN(n8626) );
  OAI211_X1 U11115 ( .C1(n8623), .C2(n8622), .A(n15003), .B(n8621), .ZN(n8624)
         );
  INV_X1 U11116 ( .A(n8624), .ZN(n8625) );
  NOR3_X1 U11117 ( .A1(n8627), .A2(n8626), .A3(n8625), .ZN(n8628) );
  OAI21_X1 U11118 ( .B1(n8849), .B2(n14993), .A(n8628), .ZN(P2_U3217) );
  OAI21_X1 U11119 ( .B1(n8629), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8630) );
  XNOR2_X1 U11120 ( .A(n8630), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10203) );
  INV_X1 U11121 ( .A(n10203), .ZN(n8889) );
  MUX2_X1 U11122 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n11907), .Z(n8829) );
  XNOR2_X1 U11123 ( .A(n8829), .B(SI_11_), .ZN(n8833) );
  INV_X1 U11124 ( .A(n10532), .ZN(n8639) );
  OAI222_X1 U11125 ( .A1(n8889), .A2(P2_U3088), .B1(n14088), .B2(n8639), .C1(
        n8633), .C2(n14086), .ZN(P2_U3316) );
  INV_X1 U11126 ( .A(n13018), .ZN(n13029) );
  OAI222_X1 U11127 ( .A1(n9579), .A2(n13618), .B1(n12508), .B2(n8634), .C1(
        n13029), .C2(P3_U3151), .ZN(P3_U3279) );
  NAND2_X1 U11128 ( .A1(n9420), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8636) );
  NAND2_X1 U11129 ( .A1(n8637), .A2(n8636), .ZN(n8827) );
  INV_X1 U11130 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8638) );
  XNOR2_X1 U11131 ( .A(n8827), .B(n8638), .ZN(n10533) );
  INV_X1 U11132 ( .A(n10533), .ZN(n9052) );
  OAI222_X1 U11133 ( .A1(n14684), .A2(n8640), .B1(P1_U3086), .B2(n9052), .C1(
        n14694), .C2(n8639), .ZN(P1_U3344) );
  INV_X1 U11134 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8649) );
  OAI211_X1 U11135 ( .C1(n8643), .C2(n8642), .A(n15003), .B(n8641), .ZN(n8648)
         );
  OAI211_X1 U11136 ( .C1(n8646), .C2(n8645), .A(n15039), .B(n8644), .ZN(n8647)
         );
  OAI211_X1 U11137 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n8649), .A(n8648), .B(
        n8647), .ZN(n8652) );
  NOR2_X1 U11138 ( .A1(n8650), .A2(n15061), .ZN(n8651) );
  AOI211_X1 U11139 ( .C1(n15052), .C2(n8653), .A(n8652), .B(n8651), .ZN(n8654)
         );
  INV_X1 U11140 ( .A(n8654), .ZN(P2_U3215) );
  INV_X1 U11141 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8655) );
  MUX2_X1 U11142 ( .A(n8655), .B(P2_REG1_REG_10__SCAN_IN), .S(n9841), .Z(n8658) );
  OAI21_X1 U11143 ( .B1(n9705), .B2(P2_REG1_REG_9__SCAN_IN), .A(n8656), .ZN(
        n8657) );
  NOR2_X1 U11144 ( .A1(n8657), .A2(n8658), .ZN(n8890) );
  AOI211_X1 U11145 ( .C1(n8658), .C2(n8657), .A(n15046), .B(n8890), .ZN(n8668)
         );
  OAI21_X1 U11146 ( .B1(n9705), .B2(P2_REG2_REG_9__SCAN_IN), .A(n8659), .ZN(
        n8662) );
  INV_X1 U11147 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8660) );
  MUX2_X1 U11148 ( .A(n8660), .B(P2_REG2_REG_10__SCAN_IN), .S(n9841), .Z(n8661) );
  INV_X1 U11149 ( .A(n15039), .ZN(n15054) );
  NOR2_X1 U11150 ( .A1(n8662), .A2(n8661), .ZN(n8884) );
  AOI211_X1 U11151 ( .C1(n8662), .C2(n8661), .A(n15054), .B(n8884), .ZN(n8667)
         );
  INV_X1 U11152 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9867) );
  NOR2_X1 U11153 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9867), .ZN(n8663) );
  AOI21_X1 U11154 ( .B1(n14987), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n8663), .ZN(
        n8664) );
  OAI21_X1 U11155 ( .B1(n8665), .B2(n14993), .A(n8664), .ZN(n8666) );
  OR3_X1 U11156 ( .A1(n8668), .A2(n8667), .A3(n8666), .ZN(P2_U3224) );
  OR2_X1 U11157 ( .A1(n8843), .A2(n8669), .ZN(n8670) );
  NAND2_X1 U11158 ( .A1(n15112), .A2(n15098), .ZN(n14015) );
  INV_X1 U11159 ( .A(n15101), .ZN(n8686) );
  NAND2_X1 U11160 ( .A1(n9834), .A2(n13563), .ZN(n9732) );
  OAI21_X1 U11161 ( .B1(n8680), .B2(n9732), .A(n8842), .ZN(n13924) );
  NAND2_X1 U11162 ( .A1(n12179), .A2(n6629), .ZN(n8673) );
  OR2_X2 U11163 ( .A1(n12498), .A2(n8673), .ZN(n13777) );
  INV_X2 U11164 ( .A(n13777), .ZN(n9326) );
  NAND2_X1 U11165 ( .A1(n12194), .A2(n12185), .ZN(n8877) );
  INV_X1 U11166 ( .A(n8877), .ZN(n8674) );
  AOI211_X1 U11167 ( .C1(n9834), .C2(n13926), .A(n6649), .B(n8674), .ZN(n13922) );
  INV_X1 U11168 ( .A(n6597), .ZN(n13808) );
  AND2_X2 U11169 ( .A1(n9117), .A2(n8675), .ZN(n13518) );
  INV_X1 U11170 ( .A(n13518), .ZN(n9357) );
  NAND2_X1 U11171 ( .A1(n6638), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8679) );
  NAND2_X1 U11172 ( .A1(n12390), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8678) );
  NAND2_X1 U11173 ( .A1(n11619), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8676) );
  INV_X1 U11174 ( .A(n13560), .ZN(n12203) );
  OAI22_X1 U11175 ( .A1(n12183), .A2(n9357), .B1(n12203), .B2(n11617), .ZN(
        n9729) );
  NAND2_X1 U11176 ( .A1(n8680), .A2(n8681), .ZN(n8683) );
  INV_X1 U11177 ( .A(n8681), .ZN(n8682) );
  NAND2_X1 U11178 ( .A1(n12447), .A2(n8682), .ZN(n8863) );
  AOI21_X1 U11179 ( .B1(n8683), .B2(n8863), .A(n13875), .ZN(n8684) );
  AOI211_X1 U11180 ( .C1(n13808), .C2(n13924), .A(n9729), .B(n8684), .ZN(
        n13929) );
  INV_X1 U11181 ( .A(n13929), .ZN(n8685) );
  AOI211_X1 U11182 ( .C1(n8686), .C2(n13924), .A(n13922), .B(n8685), .ZN(n9018) );
  MUX2_X1 U11183 ( .A(n8687), .B(n9018), .S(n15112), .Z(n8688) );
  OAI21_X1 U11184 ( .B1(n12194), .B2(n14015), .A(n8688), .ZN(P2_U3500) );
  INV_X2 U11185 ( .A(n7356), .ZN(n8696) );
  INV_X1 U11186 ( .A(n11435), .ZN(n11301) );
  INV_X1 U11187 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n8694) );
  INV_X1 U11188 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n14884) );
  OR2_X1 U11189 ( .A1(n11919), .A2(n14884), .ZN(n8699) );
  INV_X1 U11190 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8697) );
  OR2_X1 U11191 ( .A1(n9229), .A2(n8697), .ZN(n8698) );
  NAND2_X1 U11192 ( .A1(n14267), .A2(n11875), .ZN(n8709) );
  INV_X1 U11193 ( .A(n9248), .ZN(n8711) );
  NAND2_X1 U11194 ( .A1(n8711), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8708) );
  AND2_X4 U11195 ( .A1(n9248), .A2(n11935), .ZN(n11870) );
  INV_X1 U11196 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n8717) );
  NOR2_X1 U11197 ( .A1(n11907), .A2(n8705), .ZN(n8706) );
  XNOR2_X1 U11198 ( .A(n8706), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14697) );
  MUX2_X1 U11199 ( .A(n8717), .B(n14697), .S(n11404), .Z(n11936) );
  INV_X1 U11200 ( .A(n11936), .ZN(n9573) );
  NAND2_X1 U11201 ( .A1(n11870), .A2(n9573), .ZN(n8707) );
  AND3_X1 U11202 ( .A1(n8709), .A2(n8708), .A3(n8707), .ZN(n8964) );
  OR2_X2 U11203 ( .A1(n8807), .A2(n11930), .ZN(n14924) );
  AND2_X4 U11204 ( .A1(n11870), .A2(n14924), .ZN(n11874) );
  NAND2_X1 U11205 ( .A1(n11874), .A2(n14267), .ZN(n8713) );
  INV_X1 U11206 ( .A(n8967), .ZN(n8714) );
  AOI21_X1 U11207 ( .B1(n8964), .B2(n8715), .A(n8714), .ZN(n8812) );
  MUX2_X1 U11208 ( .A(n14273), .B(n8812), .S(n6663), .Z(n8718) );
  OR2_X1 U11209 ( .A1(n6663), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8716) );
  NAND2_X1 U11210 ( .A1(n9002), .A2(n8716), .ZN(n14886) );
  AND2_X1 U11211 ( .A1(n14886), .A2(n8717), .ZN(n14889) );
  AOI211_X1 U11212 ( .C1(n8718), .C2(n9002), .A(n14889), .B(n14266), .ZN(n8744) );
  XOR2_X1 U11213 ( .A(n8720), .B(n8719), .Z(n8723) );
  NAND2_X1 U11214 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n9259) );
  OAI21_X1 U11215 ( .B1(n14911), .B2(n8721), .A(n9259), .ZN(n8722) );
  AOI21_X1 U11216 ( .B1(n14901), .B2(n8723), .A(n8722), .ZN(n8730) );
  INV_X1 U11217 ( .A(n8724), .ZN(n8728) );
  NAND3_X1 U11218 ( .A1(n14289), .A2(n8726), .A3(n8725), .ZN(n8727) );
  NAND3_X1 U11219 ( .A1(n14318), .A2(n8728), .A3(n8727), .ZN(n8729) );
  OAI211_X1 U11220 ( .C1(n14320), .C2(n8731), .A(n8730), .B(n8729), .ZN(n8732)
         );
  OR2_X1 U11221 ( .A1(n8744), .A2(n8732), .ZN(P1_U3247) );
  INV_X1 U11222 ( .A(n14287), .ZN(n8733) );
  OAI211_X1 U11223 ( .C1(n8735), .C2(n8734), .A(n14318), .B(n8733), .ZN(n8742)
         );
  OAI211_X1 U11224 ( .C1(n8738), .C2(n8737), .A(n14901), .B(n8736), .ZN(n8741)
         );
  AOI22_X1 U11225 ( .A1(n14891), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n8740) );
  INV_X1 U11226 ( .A(n14320), .ZN(n14903) );
  NAND2_X1 U11227 ( .A1(n14903), .A2(n8991), .ZN(n8739) );
  NAND4_X1 U11228 ( .A1(n8742), .A2(n8741), .A3(n8740), .A4(n8739), .ZN(n8743)
         );
  OR2_X1 U11229 ( .A1(n8744), .A2(n8743), .ZN(P1_U3245) );
  INV_X1 U11230 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10386) );
  MUX2_X1 U11231 ( .A(n10386), .B(P1_REG1_REG_10__SCAN_IN), .S(n10528), .Z(
        n8747) );
  OAI21_X1 U11232 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n10380), .A(n8745), .ZN(
        n8746) );
  NOR2_X1 U11233 ( .A1(n8746), .A2(n8747), .ZN(n8817) );
  AOI211_X1 U11234 ( .C1(n8747), .C2(n8746), .A(n14323), .B(n8817), .ZN(n8758)
         );
  NAND2_X1 U11235 ( .A1(n10380), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8750) );
  INV_X1 U11236 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n8748) );
  MUX2_X1 U11237 ( .A(n8748), .B(P1_REG2_REG_10__SCAN_IN), .S(n10528), .Z(
        n8749) );
  AOI21_X1 U11238 ( .B1(n8751), .B2(n8750), .A(n8749), .ZN(n8816) );
  AND3_X1 U11239 ( .A1(n8751), .A2(n8750), .A3(n8749), .ZN(n8752) );
  NOR3_X1 U11240 ( .A1(n8816), .A2(n8752), .A3(n14906), .ZN(n8757) );
  NAND2_X1 U11241 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n14816)
         );
  INV_X1 U11242 ( .A(n14816), .ZN(n8753) );
  AOI21_X1 U11243 ( .B1(n14891), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n8753), .ZN(
        n8754) );
  OAI21_X1 U11244 ( .B1(n14320), .B2(n8755), .A(n8754), .ZN(n8756) );
  OR3_X1 U11245 ( .A1(n8758), .A2(n8757), .A3(n8756), .ZN(P1_U3253) );
  OAI222_X1 U11246 ( .A1(P3_U3151), .A2(n13044), .B1(n12508), .B2(n8759), .C1(
        n10080), .C2(n9579), .ZN(P3_U3278) );
  NAND2_X1 U11247 ( .A1(n8760), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8761) );
  MUX2_X1 U11248 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8761), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n8762) );
  AND2_X1 U11249 ( .A1(n6699), .A2(n14540), .ZN(n8764) );
  AND2_X1 U11250 ( .A1(n8805), .A2(n9249), .ZN(n12175) );
  NOR2_X1 U11251 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .ZN(
        n8768) );
  NOR4_X1 U11252 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_30__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n8767) );
  NOR4_X1 U11253 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n8766) );
  NOR4_X1 U11254 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n8765) );
  NAND4_X1 U11255 ( .A1(n8768), .A2(n8767), .A3(n8766), .A4(n8765), .ZN(n8774)
         );
  NOR4_X1 U11256 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n8772) );
  NOR4_X1 U11257 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n8771) );
  NOR4_X1 U11258 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8770) );
  NOR4_X1 U11259 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n8769) );
  NAND4_X1 U11260 ( .A1(n8772), .A2(n8771), .A3(n8770), .A4(n8769), .ZN(n8773)
         );
  OAI21_X1 U11261 ( .B1(n8774), .B2(n8773), .A(n8780), .ZN(n8802) );
  NAND2_X1 U11262 ( .A1(n14736), .A2(n11367), .ZN(n9246) );
  NAND3_X1 U11263 ( .A1(n12175), .A2(n8802), .A3(n9246), .ZN(n8777) );
  AOI21_X1 U11264 ( .B1(n8780), .B2(n8776), .A(n8775), .ZN(n8803) );
  OR2_X1 U11265 ( .A1(n8777), .A2(n8803), .ZN(n9460) );
  INV_X1 U11266 ( .A(n14986), .ZN(n14984) );
  OR2_X1 U11267 ( .A1(n14267), .A2(n11936), .ZN(n9396) );
  NAND2_X1 U11268 ( .A1(n14267), .A2(n11936), .ZN(n8782) );
  AND2_X1 U11269 ( .A1(n9396), .A2(n8782), .ZN(n12128) );
  INV_X1 U11270 ( .A(n12128), .ZN(n8796) );
  NAND2_X1 U11271 ( .A1(n8784), .A2(n14540), .ZN(n11917) );
  NOR2_X1 U11272 ( .A1(n11917), .A2(n11935), .ZN(n8783) );
  INV_X1 U11273 ( .A(n8784), .ZN(n11925) );
  NAND2_X1 U11274 ( .A1(n11925), .A2(n11367), .ZN(n11916) );
  NAND2_X1 U11275 ( .A1(n8784), .A2(n11367), .ZN(n8786) );
  OR2_X1 U11276 ( .A1(n11931), .A2(n6699), .ZN(n8785) );
  NAND2_X1 U11277 ( .A1(n14969), .A2(n14724), .ZN(n8795) );
  NAND2_X1 U11278 ( .A1(n8996), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8792) );
  INV_X1 U11279 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n8787) );
  NAND2_X1 U11280 ( .A1(n6688), .A2(n14921), .ZN(n8793) );
  OAI21_X1 U11281 ( .B1(n8807), .B2(n11936), .A(n8793), .ZN(n8794) );
  AOI21_X1 U11282 ( .B1(n8796), .B2(n8795), .A(n8794), .ZN(n14918) );
  NAND2_X1 U11283 ( .A1(n14984), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8797) );
  OAI21_X1 U11284 ( .B1(n14984), .B2(n14918), .A(n8797), .ZN(P1_U3528) );
  INV_X1 U11285 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n8801) );
  NAND2_X1 U11286 ( .A1(n15106), .A2(n8799), .ZN(n8800) );
  OAI21_X1 U11287 ( .B1(n15106), .B2(n8801), .A(n8800), .ZN(P2_U3430) );
  AND2_X1 U11288 ( .A1(n8803), .A2(n8802), .ZN(n9266) );
  NAND2_X1 U11289 ( .A1(n9266), .A2(n9459), .ZN(n9247) );
  OR2_X1 U11290 ( .A1(n9247), .A2(n8810), .ZN(n8806) );
  INV_X1 U11291 ( .A(n9246), .ZN(n8804) );
  NAND2_X1 U11292 ( .A1(n8806), .A2(n14541), .ZN(n14815) );
  INV_X1 U11293 ( .A(n14879), .ZN(n14239) );
  INV_X1 U11294 ( .A(n12175), .ZN(n9265) );
  NAND2_X1 U11295 ( .A1(n14949), .A2(n11927), .ZN(n8809) );
  NAND2_X1 U11296 ( .A1(n14815), .A2(n9249), .ZN(n9014) );
  NAND2_X1 U11297 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n9014), .ZN(n8811) );
  OAI21_X1 U11298 ( .B1(n8812), .B2(n14875), .A(n8811), .ZN(n8813) );
  AOI21_X1 U11299 ( .B1(n14217), .B2(n6688), .A(n8813), .ZN(n8814) );
  OAI21_X1 U11300 ( .B1(n11936), .B2(n14239), .A(n8814), .ZN(P1_U3232) );
  INV_X1 U11301 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n13622) );
  NAND2_X1 U11302 ( .A1(n15172), .A2(P3_U3897), .ZN(n8815) );
  OAI21_X1 U11303 ( .B1(P3_U3897), .B2(n13622), .A(n8815), .ZN(P3_U3494) );
  AOI21_X1 U11304 ( .B1(n10528), .B2(P1_REG2_REG_10__SCAN_IN), .A(n8816), .ZN(
        n9049) );
  INV_X1 U11305 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9051) );
  MUX2_X1 U11306 ( .A(n9051), .B(P1_REG2_REG_11__SCAN_IN), .S(n10533), .Z(
        n9048) );
  XNOR2_X1 U11307 ( .A(n9049), .B(n9048), .ZN(n8825) );
  AOI21_X1 U11308 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n10528), .A(n8817), .ZN(
        n8819) );
  INV_X1 U11309 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10539) );
  MUX2_X1 U11310 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10539), .S(n10533), .Z(
        n8818) );
  NAND2_X1 U11311 ( .A1(n8819), .A2(n8818), .ZN(n9055) );
  OAI21_X1 U11312 ( .B1(n8819), .B2(n8818), .A(n9055), .ZN(n8820) );
  NAND2_X1 U11313 ( .A1(n8820), .A2(n14901), .ZN(n8824) );
  NAND2_X1 U11314 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14829)
         );
  INV_X1 U11315 ( .A(n14829), .ZN(n8822) );
  NOR2_X1 U11316 ( .A1(n14320), .A2(n9052), .ZN(n8821) );
  AOI211_X1 U11317 ( .C1(n14891), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n8822), .B(
        n8821), .ZN(n8823) );
  OAI211_X1 U11318 ( .C1(n14906), .C2(n8825), .A(n8824), .B(n8823), .ZN(
        P1_U3254) );
  INV_X1 U11319 ( .A(n13058), .ZN(n13063) );
  INV_X1 U11320 ( .A(SI_18_), .ZN(n10177) );
  OAI222_X1 U11321 ( .A1(P3_U3151), .A2(n13063), .B1(n12508), .B2(n8826), .C1(
        n10177), .C2(n9579), .ZN(P3_U3277) );
  NAND2_X1 U11322 ( .A1(n8828), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9022) );
  XNOR2_X1 U11323 ( .A(n9022), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10831) );
  INV_X1 U11324 ( .A(n10831), .ZN(n9059) );
  INV_X1 U11325 ( .A(n8829), .ZN(n8831) );
  NAND2_X1 U11326 ( .A1(n8831), .A2(n8830), .ZN(n8832) );
  XNOR2_X1 U11327 ( .A(n9030), .B(SI_12_), .ZN(n9027) );
  INV_X1 U11328 ( .A(n10830), .ZN(n8839) );
  OAI222_X1 U11329 ( .A1(n9059), .A2(P1_U3086), .B1(n14684), .B2(n8835), .C1(
        n14694), .C2(n8839), .ZN(P1_U3343) );
  NAND2_X1 U11330 ( .A1(n8837), .A2(n8836), .ZN(n9546) );
  NAND2_X1 U11331 ( .A1(n9546), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8838) );
  XNOR2_X1 U11332 ( .A(n8838), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10210) );
  INV_X1 U11333 ( .A(n10210), .ZN(n9072) );
  OAI222_X1 U11334 ( .A1(P2_U3088), .A2(n9072), .B1(n14086), .B2(n8840), .C1(
        n14088), .C2(n8839), .ZN(P2_U3315) );
  INV_X1 U11335 ( .A(n13561), .ZN(n9603) );
  NAND2_X1 U11336 ( .A1(n12194), .A2(n9603), .ZN(n8841) );
  NAND2_X1 U11337 ( .A1(n8842), .A2(n8841), .ZN(n8876) );
  OR2_X1 U11339 ( .A1(n8931), .A2(n14992), .ZN(n8844) );
  INV_X1 U11340 ( .A(n12453), .ZN(n8875) );
  INV_X1 U11341 ( .A(n13916), .ZN(n9600) );
  NAND2_X1 U11342 ( .A1(n9600), .A2(n12203), .ZN(n8847) );
  NAND2_X1 U11343 ( .A1(n8874), .A2(n8847), .ZN(n8859) );
  OR2_X1 U11344 ( .A1(n8931), .A2(n8849), .ZN(n8852) );
  OR2_X1 U11345 ( .A1(n12400), .A2(n8850), .ZN(n8851) );
  OAI211_X2 U11346 ( .C1(n12399), .C2(n9217), .A(n8852), .B(n8851), .ZN(n13908) );
  NAND2_X1 U11347 ( .A1(n6638), .A2(n9097), .ZN(n8857) );
  NAND2_X1 U11348 ( .A1(n12390), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8856) );
  NAND2_X1 U11349 ( .A1(n10688), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8855) );
  NAND2_X1 U11350 ( .A1(n8853), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8854) );
  NAND4_X1 U11351 ( .A1(n8857), .A2(n8856), .A3(n8855), .A4(n8854), .ZN(n13559) );
  XNOR2_X1 U11352 ( .A(n13908), .B(n13559), .ZN(n12448) );
  INV_X1 U11353 ( .A(n12448), .ZN(n8858) );
  NAND2_X1 U11354 ( .A1(n8859), .A2(n8858), .ZN(n8930) );
  OAI21_X1 U11355 ( .B1(n8859), .B2(n8858), .A(n8930), .ZN(n13906) );
  OR2_X1 U11356 ( .A1(n8877), .A2(n13916), .ZN(n8878) );
  NAND2_X1 U11357 ( .A1(n8878), .A2(n13908), .ZN(n8860) );
  NAND2_X1 U11358 ( .A1(n8860), .A2(n9326), .ZN(n8861) );
  NOR2_X1 U11359 ( .A1(n10292), .A2(n8861), .ZN(n13907) );
  NAND2_X1 U11360 ( .A1(n9603), .A2(n13926), .ZN(n8862) );
  NAND2_X1 U11361 ( .A1(n8863), .A2(n8862), .ZN(n8880) );
  NAND2_X1 U11362 ( .A1(n8880), .A2(n12453), .ZN(n8865) );
  NAND2_X1 U11363 ( .A1(n12203), .A2(n13916), .ZN(n8864) );
  NAND2_X1 U11364 ( .A1(n8865), .A2(n8864), .ZN(n8866) );
  OAI21_X1 U11365 ( .B1(n8866), .B2(n12448), .A(n10300), .ZN(n8871) );
  NAND2_X1 U11366 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8940) );
  OAI21_X1 U11367 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n8940), .ZN(n10296) );
  INV_X1 U11368 ( .A(n10296), .ZN(n9893) );
  NAND2_X1 U11369 ( .A1(n6638), .A2(n9893), .ZN(n8870) );
  NAND2_X1 U11370 ( .A1(n12390), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8869) );
  NAND2_X1 U11371 ( .A1(n11619), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8868) );
  NAND2_X1 U11372 ( .A1(n10688), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8867) );
  NAND4_X1 U11373 ( .A1(n8870), .A2(n8869), .A3(n8868), .A4(n8867), .ZN(n13558) );
  OAI22_X1 U11374 ( .A1(n12203), .A2(n9357), .B1(n8952), .B2(n11617), .ZN(
        n9104) );
  AOI21_X1 U11375 ( .B1(n8871), .B2(n13891), .A(n9104), .ZN(n13910) );
  INV_X1 U11376 ( .A(n13910), .ZN(n8872) );
  AOI211_X1 U11377 ( .C1(n14012), .C2(n13906), .A(n13907), .B(n8872), .ZN(
        n9151) );
  AOI22_X1 U11378 ( .A1(n13992), .A2(n13908), .B1(n15109), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n8873) );
  OAI21_X1 U11379 ( .B1(n9151), .B2(n15109), .A(n8873), .ZN(P2_U3502) );
  OAI21_X1 U11380 ( .B1(n8876), .B2(n8875), .A(n8874), .ZN(n13914) );
  AOI21_X1 U11381 ( .B1(n8877), .B2(n13916), .A(n13777), .ZN(n8879) );
  AND2_X1 U11382 ( .A1(n8879), .A2(n8878), .ZN(n13915) );
  XNOR2_X1 U11383 ( .A(n8880), .B(n12453), .ZN(n8881) );
  INV_X1 U11384 ( .A(n13559), .ZN(n9889) );
  OAI22_X1 U11385 ( .A1(n9603), .A2(n9357), .B1(n9889), .B2(n11617), .ZN(n9598) );
  AOI21_X1 U11386 ( .B1(n8881), .B2(n13891), .A(n9598), .ZN(n13918) );
  INV_X1 U11387 ( .A(n13918), .ZN(n8882) );
  AOI211_X1 U11388 ( .C1(n14012), .C2(n13914), .A(n13915), .B(n8882), .ZN(
        n9364) );
  AOI22_X1 U11389 ( .A1(n13992), .A2(n13916), .B1(n15109), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n8883) );
  OAI21_X1 U11390 ( .B1(n9364), .B2(n15109), .A(n8883), .ZN(P2_U3501) );
  INV_X1 U11391 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n13661) );
  MUX2_X1 U11392 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n13661), .S(n10203), .Z(
        n8885) );
  NAND2_X1 U11393 ( .A1(n8886), .A2(n8885), .ZN(n9068) );
  OAI21_X1 U11394 ( .B1(n8886), .B2(n8885), .A(n9068), .ZN(n8896) );
  AND2_X1 U11395 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8887) );
  AOI21_X1 U11396 ( .B1(n14987), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8887), .ZN(
        n8888) );
  OAI21_X1 U11397 ( .B1(n8889), .B2(n14993), .A(n8888), .ZN(n8895) );
  INV_X1 U11398 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8891) );
  MUX2_X1 U11399 ( .A(n8891), .B(P2_REG1_REG_11__SCAN_IN), .S(n10203), .Z(
        n8892) );
  NOR2_X1 U11400 ( .A1(n8893), .A2(n8892), .ZN(n9064) );
  AOI211_X1 U11401 ( .C1(n8893), .C2(n8892), .A(n15046), .B(n9064), .ZN(n8894)
         );
  AOI211_X1 U11402 ( .C1(n15039), .C2(n8896), .A(n8895), .B(n8894), .ZN(n8897)
         );
  INV_X1 U11403 ( .A(n8897), .ZN(P2_U3225) );
  NOR2_X1 U11404 ( .A1(n8899), .A2(n8898), .ZN(n8901) );
  INV_X1 U11405 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n8900) );
  NOR2_X1 U11406 ( .A1(n8927), .A2(n8900), .ZN(P3_U3257) );
  INV_X1 U11407 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n8902) );
  NOR2_X1 U11408 ( .A1(n8927), .A2(n8902), .ZN(P3_U3236) );
  INV_X1 U11409 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n8903) );
  NOR2_X1 U11410 ( .A1(n8927), .A2(n8903), .ZN(P3_U3253) );
  INV_X1 U11411 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n8904) );
  NOR2_X1 U11412 ( .A1(n8901), .A2(n8904), .ZN(P3_U3245) );
  INV_X1 U11413 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n8905) );
  NOR2_X1 U11414 ( .A1(n8901), .A2(n8905), .ZN(P3_U3244) );
  INV_X1 U11415 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n8906) );
  NOR2_X1 U11416 ( .A1(n8901), .A2(n8906), .ZN(P3_U3243) );
  INV_X1 U11417 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n8907) );
  NOR2_X1 U11418 ( .A1(n8901), .A2(n8907), .ZN(P3_U3242) );
  INV_X1 U11419 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n8908) );
  NOR2_X1 U11420 ( .A1(n8901), .A2(n8908), .ZN(P3_U3241) );
  INV_X1 U11421 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n8909) );
  NOR2_X1 U11422 ( .A1(n8927), .A2(n8909), .ZN(P3_U3263) );
  INV_X1 U11423 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n8910) );
  NOR2_X1 U11424 ( .A1(n8901), .A2(n8910), .ZN(P3_U3262) );
  INV_X1 U11425 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n8911) );
  NOR2_X1 U11426 ( .A1(n8927), .A2(n8911), .ZN(P3_U3261) );
  INV_X1 U11427 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n8912) );
  NOR2_X1 U11428 ( .A1(n8901), .A2(n8912), .ZN(P3_U3260) );
  INV_X1 U11429 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n8913) );
  NOR2_X1 U11430 ( .A1(n8927), .A2(n8913), .ZN(P3_U3259) );
  INV_X1 U11431 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n13701) );
  NOR2_X1 U11432 ( .A1(n8901), .A2(n13701), .ZN(P3_U3258) );
  INV_X1 U11433 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n8914) );
  NOR2_X1 U11434 ( .A1(n8901), .A2(n8914), .ZN(P3_U3240) );
  INV_X1 U11435 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n8915) );
  NOR2_X1 U11436 ( .A1(n8927), .A2(n8915), .ZN(P3_U3256) );
  INV_X1 U11437 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n13687) );
  NOR2_X1 U11438 ( .A1(n8927), .A2(n13687), .ZN(P3_U3255) );
  INV_X1 U11439 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n8916) );
  NOR2_X1 U11440 ( .A1(n8927), .A2(n8916), .ZN(P3_U3254) );
  INV_X1 U11441 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n8917) );
  NOR2_X1 U11442 ( .A1(n8927), .A2(n8917), .ZN(P3_U3252) );
  INV_X1 U11443 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n8918) );
  NOR2_X1 U11444 ( .A1(n8927), .A2(n8918), .ZN(P3_U3250) );
  INV_X1 U11445 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n8919) );
  NOR2_X1 U11446 ( .A1(n8901), .A2(n8919), .ZN(P3_U3237) );
  INV_X1 U11447 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n8920) );
  NOR2_X1 U11448 ( .A1(n8901), .A2(n8920), .ZN(P3_U3238) );
  INV_X1 U11449 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n8921) );
  NOR2_X1 U11450 ( .A1(n8927), .A2(n8921), .ZN(P3_U3234) );
  INV_X1 U11451 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n8922) );
  NOR2_X1 U11452 ( .A1(n8927), .A2(n8922), .ZN(P3_U3246) );
  INV_X1 U11453 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n8923) );
  NOR2_X1 U11454 ( .A1(n8927), .A2(n8923), .ZN(P3_U3239) );
  INV_X1 U11455 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n8924) );
  NOR2_X1 U11456 ( .A1(n8927), .A2(n8924), .ZN(P3_U3249) );
  INV_X1 U11457 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n8925) );
  NOR2_X1 U11458 ( .A1(n8927), .A2(n8925), .ZN(P3_U3251) );
  INV_X1 U11459 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n13619) );
  NOR2_X1 U11460 ( .A1(n8927), .A2(n13619), .ZN(P3_U3247) );
  INV_X1 U11461 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n8926) );
  NOR2_X1 U11462 ( .A1(n8927), .A2(n8926), .ZN(P3_U3248) );
  INV_X1 U11463 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n8928) );
  NOR2_X1 U11464 ( .A1(n8927), .A2(n8928), .ZN(P3_U3235) );
  INV_X1 U11465 ( .A(n13908), .ZN(n9148) );
  NAND2_X1 U11466 ( .A1(n9148), .A2(n9889), .ZN(n8929) );
  NAND2_X1 U11467 ( .A1(n8930), .A2(n8929), .ZN(n10290) );
  NAND2_X1 U11468 ( .A1(n9238), .A2(n12393), .ZN(n8933) );
  AOI22_X1 U11469 ( .A1(n11505), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n11504), 
        .B2(n15009), .ZN(n8932) );
  NAND2_X1 U11470 ( .A1(n10290), .A2(n12451), .ZN(n10289) );
  OR2_X1 U11471 ( .A1(n15089), .A2(n13558), .ZN(n8934) );
  NAND2_X1 U11472 ( .A1(n10289), .A2(n8934), .ZN(n8948) );
  NAND2_X1 U11473 ( .A1(n9302), .A2(n12393), .ZN(n8937) );
  AOI22_X1 U11474 ( .A1(n11505), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n11504), 
        .B2(n8935), .ZN(n8936) );
  NAND2_X1 U11475 ( .A1(n8937), .A2(n8936), .ZN(n12227) );
  INV_X1 U11476 ( .A(n8940), .ZN(n8938) );
  NAND2_X1 U11477 ( .A1(n8938), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9350) );
  INV_X1 U11478 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8939) );
  NAND2_X1 U11479 ( .A1(n8940), .A2(n8939), .ZN(n8941) );
  AND2_X1 U11480 ( .A1(n9350), .A2(n8941), .ZN(n10139) );
  NAND2_X1 U11481 ( .A1(n6638), .A2(n10139), .ZN(n8946) );
  NAND2_X1 U11482 ( .A1(n12390), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8945) );
  INV_X4 U11483 ( .A(n8942), .ZN(n11619) );
  NAND2_X1 U11484 ( .A1(n11619), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8944) );
  NAND2_X1 U11485 ( .A1(n11618), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8943) );
  NAND4_X1 U11486 ( .A1(n8946), .A2(n8945), .A3(n8944), .A4(n8943), .ZN(n13557) );
  XNOR2_X1 U11487 ( .A(n12227), .B(n13557), .ZN(n12454) );
  INV_X1 U11488 ( .A(n12454), .ZN(n8947) );
  NAND2_X1 U11489 ( .A1(n8948), .A2(n8947), .ZN(n9430) );
  OAI21_X1 U11490 ( .B1(n8948), .B2(n8947), .A(n9430), .ZN(n10030) );
  INV_X1 U11491 ( .A(n15089), .ZN(n10297) );
  NAND2_X1 U11492 ( .A1(n10292), .A2(n10297), .ZN(n10293) );
  AOI21_X1 U11493 ( .B1(n10293), .B2(n12227), .A(n13777), .ZN(n8949) );
  NAND2_X1 U11494 ( .A1(n8949), .A2(n10319), .ZN(n10028) );
  INV_X1 U11495 ( .A(n10028), .ZN(n8962) );
  NAND2_X1 U11496 ( .A1(n9889), .A2(n13908), .ZN(n10299) );
  NAND2_X1 U11497 ( .A1(n10300), .A2(n10299), .ZN(n8951) );
  INV_X1 U11498 ( .A(n12451), .ZN(n8950) );
  NAND2_X1 U11499 ( .A1(n8951), .A2(n8950), .ZN(n10302) );
  NAND2_X1 U11500 ( .A1(n15089), .A2(n8952), .ZN(n8953) );
  NAND2_X1 U11501 ( .A1(n10302), .A2(n8953), .ZN(n9437) );
  XNOR2_X1 U11502 ( .A(n9437), .B(n12454), .ZN(n8960) );
  XNOR2_X1 U11503 ( .A(n9350), .B(P2_REG3_REG_6__SCAN_IN), .ZN(n9325) );
  NAND2_X1 U11504 ( .A1(n6638), .A2(n9325), .ZN(n8957) );
  NAND2_X1 U11505 ( .A1(n12390), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8956) );
  NAND2_X1 U11506 ( .A1(n11618), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8955) );
  NAND2_X1 U11507 ( .A1(n11619), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8954) );
  NAND4_X1 U11508 ( .A1(n8957), .A2(n8956), .A3(n8955), .A4(n8954), .ZN(n13556) );
  NAND2_X1 U11509 ( .A1(n13517), .A2(n13556), .ZN(n8959) );
  NAND2_X1 U11510 ( .A1(n13558), .A2(n13518), .ZN(n8958) );
  NAND2_X1 U11511 ( .A1(n8959), .A2(n8958), .ZN(n10130) );
  AOI21_X1 U11512 ( .B1(n8960), .B2(n13891), .A(n10130), .ZN(n10032) );
  INV_X1 U11513 ( .A(n10032), .ZN(n8961) );
  AOI211_X1 U11514 ( .C1(n14012), .C2(n10030), .A(n8962), .B(n8961), .ZN(n9298) );
  AOI22_X1 U11515 ( .A1(n13992), .A2(n12227), .B1(n15109), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n8963) );
  OAI21_X1 U11516 ( .B1(n9298), .B2(n15109), .A(n8963), .ZN(P2_U3504) );
  INV_X1 U11517 ( .A(n8964), .ZN(n8965) );
  NAND2_X1 U11518 ( .A1(n14265), .A2(n11875), .ZN(n8973) );
  NAND2_X1 U11519 ( .A1(n11870), .A2(n14920), .ZN(n8972) );
  NAND2_X1 U11520 ( .A1(n8973), .A2(n8972), .ZN(n8974) );
  XNOR2_X1 U11521 ( .A(n8974), .B(n11793), .ZN(n8980) );
  NAND2_X1 U11522 ( .A1(n11874), .A2(n6688), .ZN(n8977) );
  NAND2_X1 U11523 ( .A1(n11875), .A2(n14920), .ZN(n8976) );
  NAND2_X1 U11524 ( .A1(n8977), .A2(n8976), .ZN(n8978) );
  XNOR2_X1 U11525 ( .A(n8980), .B(n8978), .ZN(n9010) );
  NAND2_X1 U11526 ( .A1(n9009), .A2(n9010), .ZN(n8982) );
  INV_X1 U11527 ( .A(n8978), .ZN(n8979) );
  NAND2_X1 U11528 ( .A1(n8980), .A2(n8979), .ZN(n8981) );
  NAND2_X1 U11529 ( .A1(n11381), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8989) );
  INV_X1 U11530 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9520) );
  OR2_X1 U11531 ( .A1(n11435), .A2(n9520), .ZN(n8985) );
  OR2_X1 U11532 ( .A1(n9229), .A2(n8983), .ZN(n8984) );
  AND2_X1 U11533 ( .A1(n8985), .A2(n8984), .ZN(n8988) );
  OR2_X1 U11534 ( .A1(n11919), .A2(n8986), .ZN(n8987) );
  NAND3_X1 U11535 ( .A1(n8989), .A2(n8988), .A3(n8987), .ZN(n9387) );
  OR2_X1 U11536 ( .A1(n11391), .A2(n13734), .ZN(n8992) );
  INV_X1 U11537 ( .A(n14933), .ZN(n11945) );
  NAND2_X1 U11538 ( .A1(n6423), .A2(n11945), .ZN(n8993) );
  NAND2_X1 U11539 ( .A1(n8994), .A2(n8993), .ZN(n9212) );
  OAI22_X1 U11540 ( .A1(n11947), .A2(n8975), .B1(n14933), .B2(n11880), .ZN(
        n8995) );
  XNOR2_X1 U11541 ( .A(n8995), .B(n11793), .ZN(n9214) );
  XNOR2_X1 U11542 ( .A(n9212), .B(n9214), .ZN(n9210) );
  XOR2_X1 U11543 ( .A(n9211), .B(n9210), .Z(n9008) );
  NAND2_X1 U11544 ( .A1(n11381), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9001) );
  OR2_X1 U11545 ( .A1(n11919), .A2(n8997), .ZN(n8999) );
  OR2_X1 U11546 ( .A1(n9229), .A2(n9508), .ZN(n8998) );
  NAND4_X2 U11547 ( .A1(n9001), .A2(n9000), .A3(n8999), .A4(n8998), .ZN(n14264) );
  INV_X1 U11548 ( .A(n14264), .ZN(n9004) );
  INV_X1 U11549 ( .A(n14394), .ZN(n14517) );
  OR2_X1 U11550 ( .A1(n14233), .A2(n14517), .ZN(n14870) );
  INV_X1 U11551 ( .A(n6688), .ZN(n9576) );
  OAI22_X1 U11552 ( .A1(n9004), .A2(n14871), .B1(n14870), .B2(n9576), .ZN(
        n9006) );
  NOR2_X1 U11553 ( .A1(n14239), .A2(n14933), .ZN(n9005) );
  AOI211_X1 U11554 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n9014), .A(n9006), .B(
        n9005), .ZN(n9007) );
  OAI21_X1 U11555 ( .B1(n14875), .B2(n9008), .A(n9007), .ZN(P1_U3237) );
  XOR2_X1 U11556 ( .A(n9009), .B(n9010), .Z(n9016) );
  INV_X1 U11557 ( .A(n14267), .ZN(n9011) );
  OAI22_X1 U11558 ( .A1(n11947), .A2(n14871), .B1(n14870), .B2(n9011), .ZN(
        n9013) );
  NOR2_X1 U11559 ( .A1(n14239), .A2(n9395), .ZN(n9012) );
  AOI211_X1 U11560 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n9014), .A(n9013), .B(
        n9012), .ZN(n9015) );
  OAI21_X1 U11561 ( .B1(n14875), .B2(n9016), .A(n9015), .ZN(P1_U3222) );
  OAI222_X1 U11562 ( .A1(n12508), .A2(n9017), .B1(P3_U3151), .B2(n9776), .C1(
        n10198), .C2(n9579), .ZN(P3_U3276) );
  INV_X1 U11563 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9019) );
  MUX2_X1 U11564 ( .A(n9019), .B(n9018), .S(n15106), .Z(n9020) );
  OAI21_X1 U11565 ( .B1(n12194), .B2(n14064), .A(n9020), .ZN(P2_U3433) );
  INV_X1 U11566 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9021) );
  NAND2_X1 U11567 ( .A1(n9022), .A2(n9021), .ZN(n9023) );
  NAND2_X1 U11568 ( .A1(n9023), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9025) );
  INV_X1 U11569 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9024) );
  NAND2_X1 U11570 ( .A1(n9025), .A2(n9024), .ZN(n9081) );
  OR2_X1 U11571 ( .A1(n9025), .A2(n9024), .ZN(n9026) );
  INV_X1 U11572 ( .A(n10837), .ZN(n9645) );
  NAND2_X1 U11573 ( .A1(n9030), .A2(n9029), .ZN(n9031) );
  MUX2_X1 U11574 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n11907), .Z(n9032) );
  NAND2_X1 U11575 ( .A1(n9032), .A2(SI_13_), .ZN(n9410) );
  INV_X1 U11576 ( .A(n9032), .ZN(n9034) );
  NAND2_X1 U11577 ( .A1(n9034), .A2(n9033), .ZN(n9035) );
  NAND2_X1 U11578 ( .A1(n9410), .A2(n9035), .ZN(n9036) );
  NAND2_X1 U11579 ( .A1(n9037), .A2(n9036), .ZN(n9038) );
  AND2_X1 U11580 ( .A1(n9412), .A2(n9038), .ZN(n10836) );
  INV_X1 U11581 ( .A(n10836), .ZN(n9044) );
  OAI222_X1 U11582 ( .A1(n9645), .A2(P1_U3086), .B1(n14684), .B2(n9039), .C1(
        n14694), .C2(n9044), .ZN(P1_U3342) );
  NAND2_X1 U11583 ( .A1(n9042), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9040) );
  MUX2_X1 U11584 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9040), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n9041) );
  INV_X1 U11585 ( .A(n9041), .ZN(n9043) );
  INV_X1 U11586 ( .A(n15051), .ZN(n9046) );
  OAI222_X1 U11587 ( .A1(P2_U3088), .A2(n9046), .B1(n14086), .B2(n9045), .C1(
        n14088), .C2(n9044), .ZN(P2_U3314) );
  INV_X1 U11588 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9047) );
  AOI22_X1 U11589 ( .A1(n10831), .A2(n9047), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n9059), .ZN(n9054) );
  OR2_X1 U11590 ( .A1(n9049), .A2(n9048), .ZN(n9050) );
  OAI21_X1 U11591 ( .B1(n9052), .B2(n9051), .A(n9050), .ZN(n9053) );
  NOR2_X1 U11592 ( .A1(n9054), .A2(n9053), .ZN(n9561) );
  AOI21_X1 U11593 ( .B1(n9054), .B2(n9053), .A(n9561), .ZN(n9063) );
  INV_X1 U11594 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14750) );
  AOI22_X1 U11595 ( .A1(n10831), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n14750), 
        .B2(n9059), .ZN(n9057) );
  OAI21_X1 U11596 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n10533), .A(n9055), .ZN(
        n9056) );
  NAND2_X1 U11597 ( .A1(n9057), .A2(n9056), .ZN(n9555) );
  OAI21_X1 U11598 ( .B1(n9057), .B2(n9056), .A(n9555), .ZN(n9061) );
  AND2_X1 U11599 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n11035) );
  AOI21_X1 U11600 ( .B1(n14891), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n11035), 
        .ZN(n9058) );
  OAI21_X1 U11601 ( .B1(n14320), .B2(n9059), .A(n9058), .ZN(n9060) );
  AOI21_X1 U11602 ( .B1(n9061), .B2(n14901), .A(n9060), .ZN(n9062) );
  OAI21_X1 U11603 ( .B1(n9063), .B2(n14906), .A(n9062), .ZN(P1_U3255) );
  XOR2_X1 U11604 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n10210), .Z(n9066) );
  NAND2_X1 U11605 ( .A1(n9065), .A2(n9066), .ZN(n9900) );
  OAI21_X1 U11606 ( .B1(n9066), .B2(n9065), .A(n9900), .ZN(n9067) );
  NAND2_X1 U11607 ( .A1(n9067), .A2(n15003), .ZN(n9076) );
  INV_X1 U11608 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10366) );
  XNOR2_X1 U11609 ( .A(n10210), .B(n10366), .ZN(n9070) );
  OAI21_X1 U11610 ( .B1(n9070), .B2(n9069), .A(n9897), .ZN(n9074) );
  NAND2_X1 U11611 ( .A1(n14987), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n9071) );
  NAND2_X1 U11612 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n10228)
         );
  OAI211_X1 U11613 ( .C1(n14993), .C2(n9072), .A(n9071), .B(n10228), .ZN(n9073) );
  AOI21_X1 U11614 ( .B1(n9074), .B2(n15039), .A(n9073), .ZN(n9075) );
  NAND2_X1 U11615 ( .A1(n9076), .A2(n9075), .ZN(P2_U3226) );
  OR2_X1 U11616 ( .A1(n9407), .A2(n14068), .ZN(n9077) );
  XNOR2_X1 U11617 ( .A(n9077), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10648) );
  INV_X1 U11618 ( .A(n10648), .ZN(n10460) );
  NAND2_X1 U11619 ( .A1(n9412), .A2(n9410), .ZN(n9079) );
  XNOR2_X1 U11620 ( .A(n9409), .B(SI_14_), .ZN(n9078) );
  INV_X1 U11621 ( .A(n10968), .ZN(n9084) );
  OAI222_X1 U11622 ( .A1(n10460), .A2(P2_U3088), .B1(n14088), .B2(n9084), .C1(
        n9080), .C2(n14086), .ZN(P2_U3313) );
  NAND2_X1 U11623 ( .A1(n9081), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9082) );
  XNOR2_X1 U11624 ( .A(n9082), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10969) );
  INV_X1 U11625 ( .A(n10969), .ZN(n9651) );
  OAI222_X1 U11626 ( .A1(P1_U3086), .A2(n9651), .B1(n14694), .B2(n9084), .C1(
        n9083), .C2(n14684), .ZN(P1_U3341) );
  INV_X1 U11627 ( .A(n9087), .ZN(n9085) );
  NAND2_X1 U11628 ( .A1(n15087), .A2(n9085), .ZN(n15085) );
  OR2_X1 U11629 ( .A1(n15085), .A2(n15084), .ZN(n9086) );
  INV_X1 U11630 ( .A(n9101), .ZN(n9119) );
  INV_X1 U11631 ( .A(n12443), .ZN(n12494) );
  OR2_X1 U11632 ( .A1(n15084), .A2(n9087), .ZN(n9088) );
  OR2_X1 U11633 ( .A1(n9089), .A2(n9088), .ZN(n9090) );
  NAND2_X1 U11634 ( .A1(n9090), .A2(n9099), .ZN(n9096) );
  NOR2_X1 U11635 ( .A1(n9092), .A2(n9091), .ZN(n9094) );
  AND2_X1 U11636 ( .A1(n9094), .A2(n9093), .ZN(n9095) );
  NAND2_X1 U11637 ( .A1(n9096), .A2(n9095), .ZN(n9597) );
  AOI22_X1 U11638 ( .A1(n13495), .A2(n9097), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n9103) );
  NOR2_X1 U11639 ( .A1(n6629), .A2(n12488), .ZN(n9098) );
  NAND2_X1 U11640 ( .A1(n6667), .A2(n9098), .ZN(n9810) );
  INV_X1 U11641 ( .A(n9099), .ZN(n9100) );
  OAI21_X2 U11642 ( .B1(n9101), .B2(n9810), .A(n13825), .ZN(n13510) );
  NOR2_X1 U11643 ( .A1(n13525), .A2(n9148), .ZN(n9102) );
  AOI211_X1 U11644 ( .C1(n13521), .C2(n9104), .A(n9103), .B(n9102), .ZN(n9123)
         );
  NAND2_X1 U11645 ( .A1(n13561), .A2(n13777), .ZN(n9106) );
  NOR2_X1 U11646 ( .A1(n9732), .A2(n9326), .ZN(n9105) );
  NOR2_X1 U11647 ( .A1(n13459), .A2(n9834), .ZN(n9728) );
  NAND2_X1 U11648 ( .A1(n9602), .A2(n9106), .ZN(n9107) );
  NAND2_X1 U11649 ( .A1(n9726), .A2(n9107), .ZN(n9108) );
  XNOR2_X1 U11650 ( .A(n13459), .B(n13916), .ZN(n9109) );
  NAND2_X1 U11651 ( .A1(n13560), .A2(n13777), .ZN(n9110) );
  XNOR2_X1 U11652 ( .A(n9109), .B(n9110), .ZN(n9604) );
  INV_X1 U11653 ( .A(n9109), .ZN(n9111) );
  NAND2_X1 U11654 ( .A1(n9111), .A2(n9110), .ZN(n9112) );
  XNOR2_X1 U11655 ( .A(n13459), .B(n13908), .ZN(n9113) );
  AND2_X1 U11656 ( .A1(n13559), .A2(n13777), .ZN(n9114) );
  NAND2_X1 U11657 ( .A1(n9113), .A2(n9114), .ZN(n9327) );
  INV_X1 U11658 ( .A(n9113), .ZN(n9890) );
  INV_X1 U11659 ( .A(n9114), .ZN(n9115) );
  NAND2_X1 U11660 ( .A1(n9890), .A2(n9115), .ZN(n9116) );
  AND2_X1 U11661 ( .A1(n9327), .A2(n9116), .ZN(n9120) );
  NOR2_X1 U11662 ( .A1(n15098), .A2(n9117), .ZN(n9118) );
  NAND2_X2 U11663 ( .A1(n9119), .A2(n9118), .ZN(n13478) );
  OAI211_X1 U11664 ( .C1(n9121), .C2(n9120), .A(n13527), .B(n9329), .ZN(n9122)
         );
  NAND2_X1 U11665 ( .A1(n9123), .A2(n9122), .ZN(P2_U3190) );
  INV_X1 U11666 ( .A(n9124), .ZN(n9127) );
  NOR2_X1 U11667 ( .A1(n15085), .A2(n9125), .ZN(n9126) );
  NAND2_X1 U11668 ( .A1(n9127), .A2(n9126), .ZN(n9128) );
  NAND2_X1 U11669 ( .A1(n12489), .A2(n12441), .ZN(n9807) );
  NOR2_X1 U11670 ( .A1(n15075), .A2(n9807), .ZN(n13925) );
  INV_X1 U11671 ( .A(n13925), .ZN(n10325) );
  OAI21_X1 U11672 ( .B1(n12489), .B2(n9130), .A(n9129), .ZN(n9131) );
  INV_X1 U11673 ( .A(n13825), .ZN(n15062) );
  AOI22_X1 U11674 ( .A1(n13868), .A2(n9131), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n15062), .ZN(n9133) );
  INV_X4 U11675 ( .A(n13868), .ZN(n15075) );
  NAND2_X1 U11676 ( .A1(n15075), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9132) );
  OAI211_X1 U11677 ( .C1(n10325), .C2(n12450), .A(n9133), .B(n9132), .ZN(
        P2_U3265) );
  OR2_X1 U11678 ( .A1(n9660), .A2(P3_U3151), .ZN(n12959) );
  NAND2_X1 U11679 ( .A1(n9672), .A2(n12959), .ZN(n9144) );
  NAND2_X1 U11680 ( .A1(n9660), .A2(n12917), .ZN(n9134) );
  AND2_X1 U11681 ( .A1(n9135), .A2(n9134), .ZN(n9142) );
  MUX2_X1 U11682 ( .A(n9139), .B(P3_U3897), .S(n11665), .Z(n13071) );
  INV_X1 U11683 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n9804) );
  INV_X1 U11684 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10286) );
  MUX2_X1 U11685 ( .A(n9804), .B(n10286), .S(n13037), .Z(n9136) );
  NOR2_X1 U11686 ( .A1(n9136), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9141) );
  INV_X1 U11687 ( .A(n9137), .ZN(n9138) );
  INV_X1 U11688 ( .A(n15154), .ZN(n11139) );
  NAND2_X1 U11689 ( .A1(P3_U3897), .A2(n8044), .ZN(n13078) );
  NAND2_X1 U11690 ( .A1(n9139), .A2(n13037), .ZN(n15140) );
  NAND3_X1 U11691 ( .A1(n11139), .A2(n13078), .A3(n15140), .ZN(n9140) );
  OAI21_X1 U11692 ( .B1(n9282), .B2(n9141), .A(n9140), .ZN(n9146) );
  INV_X1 U11693 ( .A(n9142), .ZN(n9143) );
  AND2_X1 U11694 ( .A1(n9144), .A2(n9143), .ZN(n15113) );
  AOI22_X1 U11695 ( .A1(n15113), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n9145) );
  OAI211_X1 U11696 ( .C1(n15150), .C2(n9159), .A(n9146), .B(n9145), .ZN(
        P3_U3182) );
  INV_X1 U11697 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9147) );
  OAI22_X1 U11698 ( .A1(n14064), .A2(n9148), .B1(n15106), .B2(n9147), .ZN(
        n9149) );
  INV_X1 U11699 ( .A(n9149), .ZN(n9150) );
  OAI21_X1 U11700 ( .B1(n9151), .B2(n15104), .A(n9150), .ZN(P2_U3439) );
  MUX2_X1 U11701 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13037), .Z(n9365) );
  XOR2_X1 U11702 ( .A(n9190), .B(n9365), .Z(n9366) );
  INV_X1 U11703 ( .A(n9152), .ZN(n9153) );
  AOI22_X1 U11704 ( .A1(n9283), .A2(n9282), .B1(n6583), .B2(n9153), .ZN(n9193)
         );
  MUX2_X1 U11705 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n13037), .Z(n9154) );
  XOR2_X1 U11706 ( .A(n9207), .B(n9154), .Z(n9194) );
  OAI22_X1 U11707 ( .A1(n9193), .A2(n9194), .B1(n9154), .B2(n9177), .ZN(n9469)
         );
  MUX2_X1 U11708 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n13037), .Z(n9155) );
  XNOR2_X1 U11709 ( .A(n9155), .B(n9478), .ZN(n9470) );
  INV_X1 U11710 ( .A(n9155), .ZN(n9156) );
  XOR2_X1 U11711 ( .A(n9366), .B(n9367), .Z(n9192) );
  INV_X1 U11712 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n9157) );
  MUX2_X1 U11713 ( .A(n9157), .B(P3_REG1_REG_4__SCAN_IN), .S(n9190), .Z(n9168)
         );
  INV_X1 U11714 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9158) );
  MUX2_X1 U11715 ( .A(n9158), .B(P3_REG1_REG_2__SCAN_IN), .S(n9207), .Z(n9197)
         );
  AND2_X1 U11716 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n9159), .ZN(n9160) );
  OR3_X1 U11717 ( .A1(n10286), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n9162) );
  OAI21_X1 U11718 ( .B1(n9173), .B2(n9160), .A(n9162), .ZN(n9285) );
  INV_X1 U11719 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n9161) );
  NAND2_X1 U11720 ( .A1(n9197), .A2(n9196), .ZN(n9195) );
  NAND2_X1 U11721 ( .A1(n9177), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9163) );
  NAND2_X1 U11722 ( .A1(n9195), .A2(n9163), .ZN(n9164) );
  XNOR2_X1 U11723 ( .A(n9164), .B(n9478), .ZN(n9472) );
  NAND2_X1 U11724 ( .A1(n9472), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n9166) );
  NAND2_X1 U11725 ( .A1(n9164), .A2(n9179), .ZN(n9165) );
  NAND2_X1 U11726 ( .A1(n9166), .A2(n9165), .ZN(n9167) );
  NAND2_X1 U11727 ( .A1(n9167), .A2(n9168), .ZN(n9373) );
  OAI21_X1 U11728 ( .B1(n9168), .B2(n9167), .A(n9373), .ZN(n9169) );
  NAND2_X1 U11729 ( .A1(n13023), .A2(n9169), .ZN(n9188) );
  AND2_X1 U11730 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n10095) );
  AOI21_X1 U11731 ( .B1(n15113), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n10095), .ZN(
        n9187) );
  INV_X1 U11732 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n9170) );
  MUX2_X1 U11733 ( .A(n9170), .B(P3_REG2_REG_4__SCAN_IN), .S(n9190), .Z(n9184)
         );
  INV_X1 U11734 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n9171) );
  NOR2_X1 U11735 ( .A1(n9804), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9172) );
  NAND2_X1 U11736 ( .A1(n7716), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9175) );
  OAI21_X1 U11737 ( .B1(n9173), .B2(n9172), .A(n9175), .ZN(n9284) );
  INV_X1 U11738 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n9174) );
  OR2_X1 U11739 ( .A1(n9284), .A2(n9174), .ZN(n9176) );
  NAND2_X1 U11740 ( .A1(n9176), .A2(n9175), .ZN(n9200) );
  NAND2_X1 U11741 ( .A1(n9177), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9178) );
  XNOR2_X1 U11742 ( .A(n9180), .B(n9478), .ZN(n9471) );
  NAND2_X1 U11743 ( .A1(n9471), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9182) );
  NAND2_X1 U11744 ( .A1(n9180), .A2(n9179), .ZN(n9181) );
  NAND2_X1 U11745 ( .A1(n9182), .A2(n9181), .ZN(n9183) );
  NAND2_X1 U11746 ( .A1(n9183), .A2(n9184), .ZN(n9377) );
  OAI21_X1 U11747 ( .B1(n9184), .B2(n9183), .A(n9377), .ZN(n9185) );
  NAND2_X1 U11748 ( .A1(n15154), .A2(n9185), .ZN(n9186) );
  NAND3_X1 U11749 ( .A1(n9188), .A2(n9187), .A3(n9186), .ZN(n9189) );
  AOI21_X1 U11750 ( .B1(n9190), .B2(n13071), .A(n9189), .ZN(n9191) );
  OAI21_X1 U11751 ( .B1(n9192), .B2(n13078), .A(n9191), .ZN(P3_U3186) );
  XOR2_X1 U11752 ( .A(n9194), .B(n9193), .Z(n9209) );
  OAI21_X1 U11753 ( .B1(n9197), .B2(n9196), .A(n9195), .ZN(n9198) );
  NAND2_X1 U11754 ( .A1(n13023), .A2(n9198), .ZN(n9205) );
  AOI22_X1 U11755 ( .A1(n15113), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n9204) );
  OAI21_X1 U11756 ( .B1(n9201), .B2(n9200), .A(n9199), .ZN(n9202) );
  NAND2_X1 U11757 ( .A1(n15154), .A2(n9202), .ZN(n9203) );
  NAND3_X1 U11758 ( .A1(n9205), .A2(n9204), .A3(n9203), .ZN(n9206) );
  AOI21_X1 U11759 ( .B1(n9207), .B2(n13071), .A(n9206), .ZN(n9208) );
  OAI21_X1 U11760 ( .B1(n9209), .B2(n13078), .A(n9208), .ZN(P3_U3184) );
  INV_X1 U11761 ( .A(n9212), .ZN(n9213) );
  NAND2_X1 U11762 ( .A1(n9214), .A2(n9213), .ZN(n9215) );
  NAND2_X1 U11763 ( .A1(n14264), .A2(n11875), .ZN(n9222) );
  NAND2_X1 U11764 ( .A1(n11870), .A2(n14135), .ZN(n9221) );
  NAND2_X1 U11765 ( .A1(n9222), .A2(n9221), .ZN(n9223) );
  XNOR2_X1 U11766 ( .A(n9223), .B(n11881), .ZN(n9227) );
  NAND2_X1 U11767 ( .A1(n11874), .A2(n14264), .ZN(n9225) );
  NAND2_X1 U11768 ( .A1(n11825), .A2(n14135), .ZN(n9224) );
  NAND2_X1 U11769 ( .A1(n9225), .A2(n9224), .ZN(n9226) );
  NAND2_X1 U11770 ( .A1(n9227), .A2(n9226), .ZN(n9228) );
  NAND2_X1 U11771 ( .A1(n11459), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9237) );
  INV_X1 U11772 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9230) );
  INV_X1 U11773 ( .A(n9253), .ZN(n9233) );
  INV_X1 U11774 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9231) );
  INV_X1 U11775 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14136) );
  NAND2_X1 U11776 ( .A1(n9231), .A2(n14136), .ZN(n9232) );
  NAND2_X1 U11777 ( .A1(n9233), .A2(n9232), .ZN(n9401) );
  OR2_X1 U11778 ( .A1(n6575), .A2(n9401), .ZN(n9235) );
  OR2_X1 U11779 ( .A1(n11919), .A2(n9468), .ZN(n9234) );
  NAND2_X1 U11780 ( .A1(n9238), .A2(n11913), .ZN(n9240) );
  AOI22_X1 U11781 ( .A1(n11874), .A2(n14263), .B1(n11825), .B2(n11964), .ZN(
        n9241) );
  NAND2_X1 U11782 ( .A1(n9242), .A2(n9241), .ZN(n9299) );
  INV_X1 U11783 ( .A(n9299), .ZN(n9243) );
  NOR2_X1 U11784 ( .A1(n9301), .A2(n9243), .ZN(n9245) );
  INV_X1 U11785 ( .A(n14263), .ZN(n11965) );
  OAI22_X1 U11786 ( .A1(n11965), .A2(n8975), .B1(n11966), .B2(n11880), .ZN(
        n9244) );
  XNOR2_X1 U11787 ( .A(n9244), .B(n11881), .ZN(n9300) );
  XNOR2_X1 U11788 ( .A(n9245), .B(n9300), .ZN(n9264) );
  INV_X1 U11789 ( .A(n14870), .ZN(n14115) );
  AOI22_X1 U11790 ( .A1(n14879), .A2(n11964), .B1(n14115), .B2(n14264), .ZN(
        n9263) );
  NAND2_X1 U11791 ( .A1(n9247), .A2(n9246), .ZN(n9250) );
  NAND3_X1 U11792 ( .A1(n9250), .A2(n9249), .A3(n9248), .ZN(n9251) );
  NAND2_X1 U11793 ( .A1(n9251), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9252) );
  INV_X1 U11794 ( .A(n9401), .ZN(n9261) );
  NAND2_X1 U11795 ( .A1(n11381), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9258) );
  OR2_X1 U11796 ( .A1(n9229), .A2(n9688), .ZN(n9257) );
  NAND2_X1 U11797 ( .A1(n9253), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9629) );
  OAI21_X1 U11798 ( .B1(n9253), .B2(P1_REG3_REG_5__SCAN_IN), .A(n9629), .ZN(
        n9691) );
  OR2_X1 U11799 ( .A1(n11435), .A2(n9691), .ZN(n9256) );
  OR2_X1 U11800 ( .A1(n11919), .A2(n9254), .ZN(n9255) );
  INV_X1 U11801 ( .A(n14262), .ZN(n9938) );
  OAI21_X1 U11802 ( .B1(n14871), .B2(n9938), .A(n9259), .ZN(n9260) );
  AOI21_X1 U11803 ( .B1(n14236), .B2(n9261), .A(n9260), .ZN(n9262) );
  OAI211_X1 U11804 ( .C1(n9264), .C2(n14875), .A(n9263), .B(n9262), .ZN(
        P1_U3230) );
  NOR2_X1 U11805 ( .A1(n9265), .A2(n9459), .ZN(n9267) );
  NAND2_X1 U11806 ( .A1(n9267), .A2(n9266), .ZN(n11466) );
  INV_X1 U11807 ( .A(n9268), .ZN(n9269) );
  XOR2_X1 U11808 ( .A(n12131), .B(n9389), .Z(n14919) );
  AND2_X1 U11809 ( .A1(n9573), .A2(n14920), .ZN(n9270) );
  NOR2_X1 U11810 ( .A1(n9519), .A2(n9270), .ZN(n9275) );
  NOR2_X2 U11811 ( .A1(n11466), .A2(n11367), .ZN(n14739) );
  AND2_X1 U11812 ( .A1(n14739), .A2(n14736), .ZN(n11771) );
  NOR2_X1 U11813 ( .A1(n14541), .A2(n8787), .ZN(n9274) );
  INV_X1 U11814 ( .A(n9271), .ZN(n9272) );
  NAND2_X1 U11815 ( .A1(n14544), .A2(n14921), .ZN(n14525) );
  OAI22_X1 U11816 ( .A1(n9395), .A2(n14506), .B1(n14525), .B2(n11947), .ZN(
        n9273) );
  AOI211_X1 U11817 ( .C1(n9275), .C2(n11771), .A(n9274), .B(n9273), .ZN(n9281)
         );
  INV_X1 U11818 ( .A(n9275), .ZN(n14925) );
  XNOR2_X1 U11819 ( .A(n14925), .B(n9576), .ZN(n9276) );
  NOR2_X1 U11820 ( .A1(n9276), .A2(n14724), .ZN(n9279) );
  INV_X1 U11821 ( .A(n12131), .ZN(n9277) );
  AOI21_X1 U11822 ( .B1(n9277), .B2(n14267), .A(n14724), .ZN(n9278) );
  OAI22_X1 U11823 ( .A1(n9279), .A2(n14267), .B1(n9278), .B2(n14394), .ZN(
        n14923) );
  MUX2_X1 U11824 ( .A(n14923), .B(n8390), .S(n14743), .Z(n9280) );
  OAI211_X1 U11825 ( .C1(n14546), .C2(n14919), .A(n9281), .B(n9280), .ZN(
        P1_U3292) );
  XOR2_X1 U11826 ( .A(n9283), .B(n9282), .Z(n9294) );
  XNOR2_X1 U11827 ( .A(n9284), .B(P3_REG2_REG_1__SCAN_IN), .ZN(n9291) );
  AOI22_X1 U11828 ( .A1(n15113), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n9290) );
  INV_X1 U11829 ( .A(n9285), .ZN(n9287) );
  OAI21_X1 U11830 ( .B1(n9287), .B2(P3_REG1_REG_1__SCAN_IN), .A(n9286), .ZN(
        n9288) );
  NAND2_X1 U11831 ( .A1(n13023), .A2(n9288), .ZN(n9289) );
  OAI211_X1 U11832 ( .C1(n11139), .C2(n9291), .A(n9290), .B(n9289), .ZN(n9292)
         );
  AOI21_X1 U11833 ( .B1(n6583), .B2(n13071), .A(n9292), .ZN(n9293) );
  OAI21_X1 U11834 ( .B1(n13078), .B2(n9294), .A(n9293), .ZN(P3_U3183) );
  INV_X1 U11835 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9295) );
  NOR2_X1 U11836 ( .A1(n15106), .A2(n9295), .ZN(n9296) );
  AOI21_X1 U11837 ( .B1(n14051), .B2(n12227), .A(n9296), .ZN(n9297) );
  OAI21_X1 U11838 ( .B1(n9298), .B2(n15104), .A(n9297), .ZN(P2_U3445) );
  NAND2_X1 U11839 ( .A1(n9302), .A2(n11913), .ZN(n9305) );
  AOI22_X1 U11840 ( .A1(n12116), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n11366), 
        .B2(n9303), .ZN(n9304) );
  NAND2_X1 U11841 ( .A1(n9305), .A2(n9304), .ZN(n11973) );
  NAND2_X1 U11842 ( .A1(n11973), .A2(n11870), .ZN(n9307) );
  NAND2_X1 U11843 ( .A1(n14262), .A2(n11825), .ZN(n9306) );
  NAND2_X1 U11844 ( .A1(n9307), .A2(n9306), .ZN(n9308) );
  XNOR2_X1 U11845 ( .A(n9308), .B(n11793), .ZN(n9610) );
  NAND2_X1 U11846 ( .A1(n11874), .A2(n14262), .ZN(n9310) );
  NAND2_X1 U11847 ( .A1(n11973), .A2(n6423), .ZN(n9309) );
  AND2_X1 U11848 ( .A1(n9310), .A2(n9309), .ZN(n9611) );
  XNOR2_X1 U11849 ( .A(n9610), .B(n9611), .ZN(n9311) );
  XNOR2_X1 U11850 ( .A(n9615), .B(n9311), .ZN(n9324) );
  AOI22_X1 U11851 ( .A1(n14879), .A2(n11973), .B1(n14115), .B2(n14263), .ZN(
        n9323) );
  INV_X1 U11852 ( .A(n9691), .ZN(n9321) );
  NAND2_X1 U11853 ( .A1(n11459), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9318) );
  INV_X1 U11854 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9312) );
  OR2_X1 U11855 ( .A1(n11921), .A2(n9312), .ZN(n9317) );
  INV_X1 U11856 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9313) );
  XNOR2_X1 U11857 ( .A(n9629), .B(n9313), .ZN(n10011) );
  OR2_X1 U11858 ( .A1(n6575), .A2(n10011), .ZN(n9316) );
  OR2_X1 U11859 ( .A1(n11919), .A2(n9314), .ZN(n9315) );
  NAND4_X1 U11860 ( .A1(n9318), .A2(n9317), .A3(n9316), .A4(n9315), .ZN(n14261) );
  INV_X1 U11861 ( .A(n14261), .ZN(n9941) );
  OAI21_X1 U11862 ( .B1(n14871), .B2(n9941), .A(n9319), .ZN(n9320) );
  AOI21_X1 U11863 ( .B1(n14236), .B2(n9321), .A(n9320), .ZN(n9322) );
  OAI211_X1 U11864 ( .C1(n9324), .C2(n14875), .A(n9323), .B(n9322), .ZN(
        P1_U3227) );
  INV_X1 U11865 ( .A(n9325), .ZN(n10320) );
  XNOR2_X1 U11866 ( .A(n13459), .B(n15089), .ZN(n10133) );
  NAND2_X1 U11867 ( .A1(n13558), .A2(n13845), .ZN(n9330) );
  XNOR2_X1 U11868 ( .A(n10133), .B(n9330), .ZN(n9888) );
  AND2_X1 U11869 ( .A1(n9888), .A2(n9327), .ZN(n9328) );
  INV_X1 U11870 ( .A(n9330), .ZN(n9331) );
  OR2_X1 U11871 ( .A1(n10133), .A2(n9331), .ZN(n9332) );
  NAND2_X1 U11872 ( .A1(n9881), .A2(n9332), .ZN(n9333) );
  XNOR2_X1 U11873 ( .A(n12227), .B(n13459), .ZN(n9334) );
  NAND2_X1 U11874 ( .A1(n13557), .A2(n13845), .ZN(n9335) );
  XNOR2_X1 U11875 ( .A(n9334), .B(n9335), .ZN(n10134) );
  NAND2_X1 U11876 ( .A1(n9333), .A2(n10134), .ZN(n10141) );
  INV_X1 U11877 ( .A(n9334), .ZN(n9336) );
  NAND2_X1 U11878 ( .A1(n9336), .A2(n9335), .ZN(n9337) );
  NAND2_X1 U11879 ( .A1(n10141), .A2(n9337), .ZN(n9697) );
  INV_X1 U11880 ( .A(n9697), .ZN(n9346) );
  NAND2_X1 U11881 ( .A1(n9616), .A2(n12393), .ZN(n9340) );
  AOI22_X1 U11882 ( .A1(n11505), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n11504), 
        .B2(n9338), .ZN(n9339) );
  NAND2_X1 U11883 ( .A1(n9340), .A2(n9339), .ZN(n15097) );
  XNOR2_X1 U11884 ( .A(n15097), .B(n13424), .ZN(n13403) );
  NAND2_X1 U11885 ( .A1(n13556), .A2(n13845), .ZN(n9341) );
  NAND2_X1 U11886 ( .A1(n13403), .A2(n9341), .ZN(n9695) );
  INV_X1 U11887 ( .A(n9695), .ZN(n9344) );
  INV_X1 U11888 ( .A(n13403), .ZN(n9343) );
  INV_X1 U11889 ( .A(n9341), .ZN(n9342) );
  NOR2_X1 U11890 ( .A1(n9344), .A2(n9745), .ZN(n9345) );
  NAND2_X1 U11891 ( .A1(n9346), .A2(n9345), .ZN(n13406) );
  OAI211_X1 U11892 ( .C1(n9346), .C2(n9345), .A(n13406), .B(n13527), .ZN(n9362) );
  INV_X1 U11893 ( .A(n13557), .ZN(n9438) );
  INV_X1 U11894 ( .A(n9350), .ZN(n9348) );
  AND2_X1 U11895 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n9347) );
  NAND2_X1 U11896 ( .A1(n9348), .A2(n9347), .ZN(n9444) );
  INV_X1 U11897 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9349) );
  OAI21_X1 U11898 ( .B1(n9350), .B2(n9349), .A(n13710), .ZN(n9351) );
  AND2_X1 U11899 ( .A1(n9444), .A2(n9351), .ZN(n15063) );
  NAND2_X1 U11900 ( .A1(n6638), .A2(n15063), .ZN(n9356) );
  NAND2_X1 U11901 ( .A1(n12390), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9355) );
  NAND2_X1 U11902 ( .A1(n11619), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9354) );
  NAND2_X1 U11903 ( .A1(n11618), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9353) );
  NAND4_X1 U11904 ( .A1(n9356), .A2(n9355), .A3(n9354), .A4(n9353), .ZN(n13555) );
  INV_X1 U11905 ( .A(n13555), .ZN(n9750) );
  OAI22_X1 U11906 ( .A1(n9438), .A2(n9357), .B1(n9750), .B2(n11617), .ZN(
        n10315) );
  INV_X1 U11907 ( .A(n10315), .ZN(n9359) );
  OAI21_X1 U11908 ( .B1(n13503), .B2(n9359), .A(n9358), .ZN(n9360) );
  AOI21_X1 U11909 ( .B1(n15097), .B2(n13510), .A(n9360), .ZN(n9361) );
  OAI211_X1 U11910 ( .C1(n13495), .C2(n10320), .A(n9362), .B(n9361), .ZN(
        P2_U3211) );
  AOI22_X1 U11911 ( .A1(n14051), .A2(n13916), .B1(n15104), .B2(
        P2_REG0_REG_2__SCAN_IN), .ZN(n9363) );
  OAI21_X1 U11912 ( .B1(n9364), .B2(n15104), .A(n9363), .ZN(P2_U3436) );
  INV_X1 U11913 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n9368) );
  INV_X1 U11914 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n9374) );
  MUX2_X1 U11915 ( .A(n9368), .B(n9374), .S(n13037), .Z(n9369) );
  NAND2_X1 U11916 ( .A1(n9369), .A2(n9384), .ZN(n15122) );
  MUX2_X1 U11917 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n13037), .Z(n9370) );
  NAND2_X1 U11918 ( .A1(n9370), .A2(n9967), .ZN(n9975) );
  NAND2_X1 U11919 ( .A1(n15122), .A2(n9975), .ZN(n9371) );
  XNOR2_X1 U11920 ( .A(n9976), .B(n9371), .ZN(n9386) );
  NAND2_X1 U11921 ( .A1(n9375), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9372) );
  NAND2_X1 U11922 ( .A1(n9373), .A2(n9372), .ZN(n9966) );
  XNOR2_X1 U11923 ( .A(n9966), .B(n9384), .ZN(n9968) );
  XNOR2_X1 U11924 ( .A(n9968), .B(n9374), .ZN(n9382) );
  NAND2_X1 U11925 ( .A1(n9375), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9376) );
  NAND2_X1 U11926 ( .A1(n9377), .A2(n9376), .ZN(n9960) );
  XNOR2_X1 U11927 ( .A(n9960), .B(n9384), .ZN(n9961) );
  XNOR2_X1 U11928 ( .A(n9961), .B(P3_REG2_REG_5__SCAN_IN), .ZN(n9378) );
  NAND2_X1 U11929 ( .A1(n15154), .A2(n9378), .ZN(n9381) );
  NOR2_X1 U11930 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9379), .ZN(n10264) );
  AOI21_X1 U11931 ( .B1(n15113), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n10264), .ZN(
        n9380) );
  OAI211_X1 U11932 ( .C1(n9382), .C2(n15140), .A(n9381), .B(n9380), .ZN(n9383)
         );
  AOI21_X1 U11933 ( .B1(n9384), .B2(n13071), .A(n9383), .ZN(n9385) );
  OAI21_X1 U11934 ( .B1(n9386), .B2(n13078), .A(n9385), .ZN(P3_U3187) );
  AND2_X1 U11935 ( .A1(n9387), .A2(n14933), .ZN(n11952) );
  OR2_X2 U11936 ( .A1(n9387), .A2(n14933), .ZN(n11956) );
  NAND2_X1 U11937 ( .A1(n11947), .A2(n14933), .ZN(n9391) );
  NAND2_X1 U11938 ( .A1(n9392), .A2(n9391), .ZN(n9502) );
  NAND2_X1 U11939 ( .A1(n14264), .A2(n14938), .ZN(n11954) );
  OR2_X1 U11940 ( .A1(n14264), .A2(n14135), .ZN(n9393) );
  OR2_X1 U11941 ( .A1(n14263), .A2(n11964), .ZN(n9678) );
  NAND2_X1 U11942 ( .A1(n14263), .A2(n11964), .ZN(n9681) );
  NAND2_X1 U11943 ( .A1(n9678), .A2(n9681), .ZN(n12127) );
  XNOR2_X1 U11944 ( .A(n9680), .B(n12127), .ZN(n9464) );
  INV_X1 U11945 ( .A(n9516), .ZN(n12130) );
  OR2_X1 U11946 ( .A1(n6688), .A2(n9395), .ZN(n9397) );
  NAND2_X1 U11947 ( .A1(n12130), .A2(n9522), .ZN(n9503) );
  NAND2_X1 U11948 ( .A1(n9503), .A2(n11956), .ZN(n9398) );
  NAND2_X1 U11949 ( .A1(n9398), .A2(n12129), .ZN(n9506) );
  NAND2_X1 U11950 ( .A1(n9506), .A2(n11957), .ZN(n9683) );
  XNOR2_X1 U11951 ( .A(n9683), .B(n12127), .ZN(n9399) );
  AOI222_X1 U11952 ( .A1(n14832), .A2(n9399), .B1(n14262), .B2(n14921), .C1(
        n14264), .C2(n14394), .ZN(n9463) );
  MUX2_X1 U11953 ( .A(n8391), .B(n9463), .S(n14544), .Z(n9405) );
  INV_X1 U11954 ( .A(n11771), .ZN(n10553) );
  NAND2_X1 U11955 ( .A1(n9519), .A2(n14933), .ZN(n9518) );
  NAND2_X1 U11956 ( .A1(n9509), .A2(n11966), .ZN(n9690) );
  OR2_X1 U11957 ( .A1(n9509), .A2(n11966), .ZN(n9400) );
  AND2_X1 U11958 ( .A1(n9690), .A2(n9400), .ZN(n9461) );
  INV_X1 U11959 ( .A(n9461), .ZN(n9402) );
  OAI22_X1 U11960 ( .A1(n10553), .A2(n9402), .B1(n9401), .B2(n14541), .ZN(
        n9403) );
  AOI21_X1 U11961 ( .B1(n14733), .B2(n11964), .A(n9403), .ZN(n9404) );
  OAI211_X1 U11962 ( .C1(n9464), .C2(n14546), .A(n9405), .B(n9404), .ZN(
        P1_U3289) );
  NAND2_X1 U11963 ( .A1(n9407), .A2(n9406), .ZN(n9542) );
  NAND2_X1 U11964 ( .A1(n9542), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9408) );
  XNOR2_X1 U11965 ( .A(n9408), .B(P2_IR_REG_15__SCAN_IN), .ZN(n10682) );
  INV_X1 U11966 ( .A(n10682), .ZN(n10623) );
  OAI21_X1 U11967 ( .B1(n9414), .B2(n9413), .A(n9410), .ZN(n9411) );
  MUX2_X1 U11968 ( .A(n9428), .B(n9415), .S(n11907), .Z(n9539) );
  XNOR2_X1 U11969 ( .A(n9539), .B(SI_15_), .ZN(n9536) );
  XNOR2_X1 U11970 ( .A(n9537), .B(n9536), .ZN(n11178) );
  INV_X1 U11971 ( .A(n11178), .ZN(n9427) );
  OAI222_X1 U11972 ( .A1(P2_U3088), .A2(n10623), .B1(n14086), .B2(n9415), .C1(
        n14088), .C2(n9427), .ZN(P2_U3312) );
  INV_X1 U11973 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9418) );
  NAND4_X1 U11974 ( .A1(n9416), .A2(n9419), .A3(n9418), .A4(n9417), .ZN(n9421)
         );
  NOR2_X1 U11975 ( .A1(n9421), .A2(n9420), .ZN(n9423) );
  NAND2_X1 U11976 ( .A1(n9423), .A2(n9422), .ZN(n9425) );
  NAND2_X1 U11977 ( .A1(n9425), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9424) );
  MUX2_X1 U11978 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9424), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n9426) );
  INV_X1 U11979 ( .A(n14902), .ZN(n10481) );
  OAI222_X1 U11980 ( .A1(n10481), .A2(P1_U3086), .B1(n14684), .B2(n9428), .C1(
        n14694), .C2(n9427), .ZN(P1_U3340) );
  OR2_X1 U11981 ( .A1(n12227), .A2(n13557), .ZN(n9429) );
  NAND2_X1 U11982 ( .A1(n9430), .A2(n9429), .ZN(n10309) );
  XNOR2_X1 U11983 ( .A(n15097), .B(n13556), .ZN(n12456) );
  NAND2_X1 U11984 ( .A1(n10309), .A2(n7209), .ZN(n10308) );
  OR2_X1 U11985 ( .A1(n15097), .A2(n13556), .ZN(n9431) );
  NAND2_X1 U11986 ( .A1(n10308), .A2(n9431), .ZN(n9435) );
  OR2_X1 U11987 ( .A1(n9925), .A2(n12399), .ZN(n9434) );
  AOI22_X1 U11988 ( .A1(n11505), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n11504), 
        .B2(n9432), .ZN(n9433) );
  XNOR2_X1 U11989 ( .A(n13414), .B(n9750), .ZN(n12458) );
  OAI21_X1 U11990 ( .B1(n9435), .B2(n12458), .A(n9482), .ZN(n15071) );
  INV_X1 U11991 ( .A(n10318), .ZN(n9436) );
  INV_X1 U11992 ( .A(n13414), .ZN(n15068) );
  AOI211_X1 U11993 ( .C1(n13414), .C2(n9436), .A(n6649), .B(n9498), .ZN(n15065) );
  NAND2_X1 U11994 ( .A1(n9437), .A2(n12454), .ZN(n9440) );
  NAND2_X1 U11995 ( .A1(n12227), .A2(n9438), .ZN(n9439) );
  NAND2_X1 U11996 ( .A1(n9440), .A2(n9439), .ZN(n10312) );
  INV_X1 U11997 ( .A(n13556), .ZN(n13404) );
  NAND2_X1 U11998 ( .A1(n15097), .A2(n13404), .ZN(n9441) );
  XOR2_X1 U11999 ( .A(n12458), .B(n9485), .Z(n9452) );
  INV_X1 U12000 ( .A(n9444), .ZN(n9442) );
  NAND2_X1 U12001 ( .A1(n9442), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9489) );
  INV_X1 U12002 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9443) );
  NAND2_X1 U12003 ( .A1(n9444), .A2(n9443), .ZN(n9445) );
  AND2_X1 U12004 ( .A1(n9489), .A2(n9445), .ZN(n9996) );
  NAND2_X1 U12005 ( .A1(n6638), .A2(n9996), .ZN(n9449) );
  NAND2_X1 U12006 ( .A1(n12390), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9448) );
  NAND2_X1 U12007 ( .A1(n11619), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9447) );
  NAND2_X1 U12008 ( .A1(n11618), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9446) );
  NAND4_X1 U12009 ( .A1(n9449), .A2(n9448), .A3(n9447), .A4(n9446), .ZN(n13554) );
  NAND2_X1 U12010 ( .A1(n13517), .A2(n13554), .ZN(n9451) );
  NAND2_X1 U12011 ( .A1(n13556), .A2(n13518), .ZN(n9450) );
  NAND2_X1 U12012 ( .A1(n9451), .A2(n9450), .ZN(n13411) );
  AOI21_X1 U12013 ( .B1(n9452), .B2(n13891), .A(n13411), .ZN(n15074) );
  INV_X1 U12014 ( .A(n15074), .ZN(n9453) );
  AOI211_X1 U12015 ( .C1(n14012), .C2(n15071), .A(n15065), .B(n9453), .ZN(
        n9458) );
  INV_X1 U12016 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9454) );
  OAI22_X1 U12017 ( .A1(n14064), .A2(n15068), .B1(n15106), .B2(n9454), .ZN(
        n9455) );
  INV_X1 U12018 ( .A(n9455), .ZN(n9456) );
  OAI21_X1 U12019 ( .B1(n9458), .B2(n15104), .A(n9456), .ZN(P2_U3451) );
  AOI22_X1 U12020 ( .A1(n13992), .A2(n13414), .B1(n15109), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n9457) );
  OAI21_X1 U12021 ( .B1(n9458), .B2(n15109), .A(n9457), .ZN(P2_U3506) );
  AOI22_X1 U12022 ( .A1(n9461), .A2(n14736), .B1(n11964), .B2(n14961), .ZN(
        n9462) );
  OAI211_X1 U12023 ( .C1(n14969), .C2(n9464), .A(n9463), .B(n9462), .ZN(n9466)
         );
  NAND2_X1 U12024 ( .A1(n9466), .A2(n14953), .ZN(n9465) );
  OAI21_X1 U12025 ( .B1(n14953), .B2(n9230), .A(n9465), .ZN(P1_U3471) );
  NAND2_X1 U12026 ( .A1(n9466), .A2(n14986), .ZN(n9467) );
  OAI21_X1 U12027 ( .B1(n14986), .B2(n9468), .A(n9467), .ZN(P1_U3532) );
  XOR2_X1 U12028 ( .A(n9470), .B(n9469), .Z(n9480) );
  INV_X1 U12029 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10051) );
  XNOR2_X1 U12030 ( .A(n9471), .B(n10051), .ZN(n9476) );
  NOR2_X1 U12031 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7724), .ZN(n10064) );
  XOR2_X1 U12032 ( .A(n9472), .B(P3_REG1_REG_3__SCAN_IN), .Z(n9473) );
  NOR2_X1 U12033 ( .A1(n15140), .A2(n9473), .ZN(n9474) );
  AOI211_X1 U12034 ( .C1(n15113), .C2(P3_ADDR_REG_3__SCAN_IN), .A(n10064), .B(
        n9474), .ZN(n9475) );
  OAI21_X1 U12035 ( .B1(n9476), .B2(n11139), .A(n9475), .ZN(n9477) );
  AOI21_X1 U12036 ( .B1(n9478), .B2(n13071), .A(n9477), .ZN(n9479) );
  OAI21_X1 U12037 ( .B1(n9480), .B2(n13078), .A(n9479), .ZN(P3_U3185) );
  NAND2_X1 U12038 ( .A1(n15068), .A2(n9750), .ZN(n9481) );
  AOI22_X1 U12039 ( .A1(n11505), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n11504), 
        .B2(n9483), .ZN(n9484) );
  XNOR2_X1 U12040 ( .A(n12245), .B(n13554), .ZN(n12459) );
  INV_X1 U12041 ( .A(n12459), .ZN(n9486) );
  OAI21_X1 U12042 ( .B1(n6552), .B2(n9486), .A(n9760), .ZN(n9999) );
  AOI21_X1 U12043 ( .B1(n9487), .B2(n9486), .A(n13875), .ZN(n9497) );
  OR2_X2 U12044 ( .A1(n9487), .A2(n9486), .ZN(n9765) );
  NAND2_X1 U12045 ( .A1(n9489), .A2(n9488), .ZN(n9490) );
  AND2_X1 U12046 ( .A1(n9709), .A2(n9490), .ZN(n9811) );
  NAND2_X1 U12047 ( .A1(n6638), .A2(n9811), .ZN(n9494) );
  NAND2_X1 U12048 ( .A1(n12390), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n9493) );
  NAND2_X1 U12049 ( .A1(n11619), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9492) );
  NAND2_X1 U12050 ( .A1(n11618), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9491) );
  NAND4_X1 U12051 ( .A1(n9494), .A2(n9493), .A3(n9492), .A4(n9491), .ZN(n13553) );
  NAND2_X1 U12052 ( .A1(n13517), .A2(n13553), .ZN(n9496) );
  NAND2_X1 U12053 ( .A1(n13555), .A2(n13518), .ZN(n9495) );
  NAND2_X1 U12054 ( .A1(n9496), .A2(n9495), .ZN(n9752) );
  AOI21_X1 U12055 ( .B1(n9497), .B2(n9765), .A(n9752), .ZN(n10004) );
  INV_X1 U12056 ( .A(n12245), .ZN(n9754) );
  NAND2_X1 U12057 ( .A1(n9498), .A2(n9754), .ZN(n9761) );
  OAI211_X1 U12058 ( .C1(n9498), .C2(n9754), .A(n9326), .B(n9761), .ZN(n9995)
         );
  OAI211_X1 U12059 ( .C1(n9999), .C2(n15093), .A(n10004), .B(n9995), .ZN(n9551) );
  INV_X1 U12060 ( .A(n9551), .ZN(n9500) );
  AOI22_X1 U12061 ( .A1(n13992), .A2(n12245), .B1(n15109), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n9499) );
  OAI21_X1 U12062 ( .B1(n9500), .B2(n15109), .A(n9499), .ZN(P2_U3507) );
  OAI222_X1 U12063 ( .A1(n9579), .A2(n10185), .B1(P3_U3151), .B2(n9775), .C1(
        n12508), .C2(n9501), .ZN(P3_U3275) );
  XNOR2_X1 U12064 ( .A(n9502), .B(n9504), .ZN(n14942) );
  INV_X1 U12065 ( .A(n14942), .ZN(n9515) );
  OR2_X1 U12066 ( .A1(n11935), .A2(n14540), .ZN(n11928) );
  OAI22_X1 U12067 ( .A1(n11965), .A2(n14637), .B1(n11947), .B2(n14517), .ZN(
        n14134) );
  NAND3_X1 U12068 ( .A1(n9503), .A2(n11956), .A3(n9504), .ZN(n9505) );
  AOI21_X1 U12069 ( .B1(n9506), .B2(n9505), .A(n14724), .ZN(n9507) );
  AOI211_X1 U12070 ( .C1(n14729), .C2(n14942), .A(n14134), .B(n9507), .ZN(
        n14939) );
  MUX2_X1 U12071 ( .A(n9508), .B(n14939), .S(n14544), .Z(n9514) );
  INV_X1 U12072 ( .A(n9518), .ZN(n9511) );
  INV_X1 U12073 ( .A(n9509), .ZN(n9510) );
  OAI211_X1 U12074 ( .C1(n14938), .C2(n9511), .A(n9510), .B(n14736), .ZN(
        n14937) );
  OAI22_X1 U12075 ( .A1(n14486), .A2(n14937), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14541), .ZN(n9512) );
  AOI21_X1 U12076 ( .B1(n14733), .B2(n14135), .A(n9512), .ZN(n9513) );
  OAI211_X1 U12077 ( .C1(n9515), .C2(n14508), .A(n9514), .B(n9513), .ZN(
        P1_U3290) );
  XNOR2_X1 U12078 ( .A(n9517), .B(n9516), .ZN(n14930) );
  INV_X1 U12079 ( .A(n14930), .ZN(n9532) );
  OAI211_X1 U12080 ( .C1(n9519), .C2(n14933), .A(n14736), .B(n9518), .ZN(
        n14931) );
  OAI22_X1 U12081 ( .A1(n14486), .A2(n14931), .B1(n9520), .B2(n14541), .ZN(
        n9521) );
  AOI21_X1 U12082 ( .B1(n14733), .B2(n11945), .A(n9521), .ZN(n9531) );
  NAND2_X1 U12083 ( .A1(n14930), .A2(n14729), .ZN(n9528) );
  OAI21_X1 U12084 ( .B1(n12130), .B2(n9522), .A(n9503), .ZN(n9526) );
  NAND2_X1 U12085 ( .A1(n6688), .A2(n14394), .ZN(n9524) );
  NAND2_X1 U12086 ( .A1(n14264), .A2(n14921), .ZN(n9523) );
  NAND2_X1 U12087 ( .A1(n9524), .A2(n9523), .ZN(n9525) );
  AOI21_X1 U12088 ( .B1(n9526), .B2(n14832), .A(n9525), .ZN(n9527) );
  NAND2_X1 U12089 ( .A1(n9528), .A2(n9527), .ZN(n14934) );
  MUX2_X1 U12090 ( .A(n14934), .B(P1_REG2_REG_2__SCAN_IN), .S(n14743), .Z(
        n9529) );
  INV_X1 U12091 ( .A(n9529), .ZN(n9530) );
  OAI211_X1 U12092 ( .C1(n9532), .C2(n14508), .A(n9531), .B(n9530), .ZN(
        P1_U3291) );
  NAND2_X1 U12093 ( .A1(n9534), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9533) );
  MUX2_X1 U12094 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9533), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n9535) );
  NAND2_X1 U12095 ( .A1(n9535), .A2(n10084), .ZN(n11054) );
  NAND2_X1 U12096 ( .A1(n9539), .A2(n9538), .ZN(n9540) );
  MUX2_X1 U12097 ( .A(n9541), .B(n13726), .S(n11907), .Z(n9585) );
  XNOR2_X1 U12098 ( .A(n9585), .B(SI_16_), .ZN(n9583) );
  XNOR2_X1 U12099 ( .A(n9584), .B(n9583), .ZN(n11168) );
  INV_X1 U12100 ( .A(n11168), .ZN(n9548) );
  OAI222_X1 U12101 ( .A1(n11054), .A2(P1_U3086), .B1(n14684), .B2(n9541), .C1(
        n14694), .C2(n9548), .ZN(P1_U3339) );
  OAI21_X1 U12102 ( .B1(n9542), .B2(P2_IR_REG_15__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9543) );
  MUX2_X1 U12103 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9543), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n9547) );
  INV_X1 U12104 ( .A(n9544), .ZN(n9545) );
  OR2_X1 U12105 ( .A1(n9546), .A2(n9545), .ZN(n9589) );
  AND2_X1 U12106 ( .A1(n9547), .A2(n9589), .ZN(n10923) );
  INV_X1 U12107 ( .A(n10923), .ZN(n10638) );
  OAI222_X1 U12108 ( .A1(P2_U3088), .A2(n10638), .B1(n14086), .B2(n13726), 
        .C1(n14088), .C2(n9548), .ZN(P2_U3311) );
  INV_X1 U12109 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9549) );
  OAI22_X1 U12110 ( .A1(n14064), .A2(n9754), .B1(n15106), .B2(n9549), .ZN(
        n9550) );
  AOI21_X1 U12111 ( .B1(n9551), .B2(n15106), .A(n9550), .ZN(n9552) );
  INV_X1 U12112 ( .A(n9552), .ZN(P2_U3454) );
  NAND2_X1 U12113 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n11216)
         );
  INV_X1 U12114 ( .A(n11216), .ZN(n9553) );
  AOI21_X1 U12115 ( .B1(n14891), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n9553), .ZN(
        n9554) );
  INV_X1 U12116 ( .A(n9554), .ZN(n9559) );
  OAI21_X1 U12117 ( .B1(n10831), .B2(P1_REG1_REG_12__SCAN_IN), .A(n9555), .ZN(
        n9557) );
  INV_X1 U12118 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10843) );
  MUX2_X1 U12119 ( .A(n10843), .B(P1_REG1_REG_13__SCAN_IN), .S(n10837), .Z(
        n9556) );
  NOR2_X1 U12120 ( .A1(n9556), .A2(n9557), .ZN(n9641) );
  AOI211_X1 U12121 ( .C1(n9557), .C2(n9556), .A(n9641), .B(n14323), .ZN(n9558)
         );
  AOI211_X1 U12122 ( .C1(n14903), .C2(n10837), .A(n9559), .B(n9558), .ZN(n9565) );
  NOR2_X1 U12123 ( .A1(n10831), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9560) );
  NOR2_X1 U12124 ( .A1(n9561), .A2(n9560), .ZN(n9563) );
  INV_X1 U12125 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10855) );
  MUX2_X1 U12126 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n10855), .S(n10837), .Z(
        n9562) );
  NAND2_X1 U12127 ( .A1(n9562), .A2(n9563), .ZN(n9644) );
  OAI211_X1 U12128 ( .C1(n9563), .C2(n9562), .A(n14318), .B(n9644), .ZN(n9564)
         );
  NAND2_X1 U12129 ( .A1(n9565), .A2(n9564), .ZN(P1_U3256) );
  NAND2_X1 U12130 ( .A1(n15193), .A2(n12771), .ZN(n12768) );
  INV_X1 U12131 ( .A(n12768), .ZN(n9566) );
  NOR2_X1 U12132 ( .A1(n15190), .A2(n9566), .ZN(n12930) );
  INV_X1 U12133 ( .A(n9665), .ZN(n9567) );
  NAND2_X1 U12134 ( .A1(n9567), .A2(n15226), .ZN(n9656) );
  AND2_X1 U12135 ( .A1(n15198), .A2(n9656), .ZN(n9568) );
  OR2_X1 U12136 ( .A1(n12930), .A2(n9568), .ZN(n9570) );
  OR2_X1 U12137 ( .A1(n9780), .A2(n14776), .ZN(n9569) );
  AND2_X1 U12138 ( .A1(n9570), .A2(n9569), .ZN(n10287) );
  INV_X1 U12139 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n9571) );
  MUX2_X1 U12140 ( .A(n10287), .B(n9571), .S(n15234), .Z(n9572) );
  OAI21_X1 U12141 ( .B1(n12771), .B2(n13384), .A(n9572), .ZN(P3_U3390) );
  OAI21_X1 U12142 ( .B1(n14733), .B2(n11771), .A(n9573), .ZN(n9575) );
  INV_X1 U12143 ( .A(n14541), .ZN(n14732) );
  AOI22_X1 U12144 ( .A1(n14743), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n14732), .ZN(n9574) );
  OAI211_X1 U12145 ( .C1(n9576), .C2(n14525), .A(n9575), .B(n9574), .ZN(n9578)
         );
  INV_X1 U12146 ( .A(n14480), .ZN(n14476) );
  AOI21_X1 U12147 ( .B1(n14476), .B2(n14546), .A(n12128), .ZN(n9577) );
  OR2_X1 U12148 ( .A1(n9578), .A2(n9577), .ZN(P1_U3293) );
  INV_X1 U12149 ( .A(SI_21_), .ZN(n9580) );
  OAI222_X1 U12150 ( .A1(P3_U3151), .A2(n10042), .B1(n12508), .B2(n9581), .C1(
        n9580), .C2(n9579), .ZN(P3_U3274) );
  NAND2_X1 U12151 ( .A1(n10084), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9582) );
  XNOR2_X1 U12152 ( .A(n9582), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14295) );
  INV_X1 U12153 ( .A(n14295), .ZN(n14300) );
  NAND2_X1 U12154 ( .A1(n9584), .A2(n9583), .ZN(n9587) );
  NAND2_X1 U12155 ( .A1(n9585), .A2(n13618), .ZN(n9586) );
  XNOR2_X1 U12156 ( .A(n10078), .B(n10077), .ZN(n11353) );
  INV_X1 U12157 ( .A(n11353), .ZN(n9595) );
  OAI222_X1 U12158 ( .A1(n14300), .A2(P1_U3086), .B1(n14689), .B2(n9588), .C1(
        n14694), .C2(n9595), .ZN(P1_U3338) );
  NAND2_X1 U12159 ( .A1(n9589), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9590) );
  MUX2_X1 U12160 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9590), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n9591) );
  INV_X1 U12161 ( .A(n9591), .ZN(n9594) );
  NOR2_X1 U12162 ( .A1(n9594), .A2(n9593), .ZN(n11256) );
  INV_X1 U12163 ( .A(n11256), .ZN(n10908) );
  OAI222_X1 U12164 ( .A1(P2_U3088), .A2(n10908), .B1(n14086), .B2(n9596), .C1(
        n14088), .C2(n9595), .ZN(P2_U3310) );
  OR2_X1 U12165 ( .A1(n9597), .A2(P2_U3088), .ZN(n9837) );
  INV_X1 U12166 ( .A(n9598), .ZN(n9599) );
  OAI22_X1 U12167 ( .A1(n13525), .A2(n9600), .B1(n9599), .B2(n13503), .ZN(
        n9601) );
  AOI21_X1 U12168 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n9837), .A(n9601), .ZN(
        n9608) );
  OAI22_X1 U12169 ( .A1(n13512), .A2(n9603), .B1(n9602), .B2(n13478), .ZN(
        n9606) );
  INV_X1 U12170 ( .A(n9604), .ZN(n9605) );
  NAND3_X1 U12171 ( .A1(n9606), .A2(n9605), .A3(n9726), .ZN(n9607) );
  OAI211_X1 U12172 ( .C1(n13478), .C2(n9609), .A(n9608), .B(n9607), .ZN(
        P2_U3209) );
  INV_X1 U12173 ( .A(n9610), .ZN(n9613) );
  INV_X1 U12174 ( .A(n9611), .ZN(n9612) );
  NAND2_X1 U12175 ( .A1(n9613), .A2(n9612), .ZN(n9614) );
  NAND2_X1 U12176 ( .A1(n9616), .A2(n11913), .ZN(n9619) );
  AOI22_X1 U12177 ( .A1(n12116), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11366), 
        .B2(n9617), .ZN(n9618) );
  NAND2_X1 U12178 ( .A1(n9619), .A2(n9618), .ZN(n14944) );
  NAND2_X1 U12179 ( .A1(n14944), .A2(n11870), .ZN(n9621) );
  NAND2_X1 U12180 ( .A1(n14261), .A2(n11825), .ZN(n9620) );
  NAND2_X1 U12181 ( .A1(n9621), .A2(n9620), .ZN(n9622) );
  XNOR2_X1 U12182 ( .A(n9622), .B(n11793), .ZN(n9624) );
  AOI22_X1 U12183 ( .A1(n14944), .A2(n11825), .B1(n11874), .B2(n14261), .ZN(
        n9623) );
  OR2_X1 U12184 ( .A1(n9624), .A2(n9623), .ZN(n10109) );
  NAND2_X1 U12185 ( .A1(n6558), .A2(n10109), .ZN(n9625) );
  XNOR2_X1 U12186 ( .A(n10110), .B(n9625), .ZN(n9640) );
  AOI22_X1 U12187 ( .A1(n14879), .A2(n14944), .B1(n14115), .B2(n14262), .ZN(
        n9639) );
  NAND2_X1 U12188 ( .A1(n11459), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9635) );
  INV_X1 U12189 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9626) );
  OR2_X1 U12190 ( .A1(n11921), .A2(n9626), .ZN(n9634) );
  INV_X1 U12191 ( .A(n9629), .ZN(n9627) );
  AOI21_X1 U12192 ( .B1(n9627), .B2(P1_REG3_REG_6__SCAN_IN), .A(
        P1_REG3_REG_7__SCAN_IN), .ZN(n9630) );
  NAND2_X1 U12193 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n9628) );
  NOR2_X1 U12194 ( .A1(n9629), .A2(n9628), .ZN(n9931) );
  OR2_X1 U12195 ( .A1(n9630), .A2(n9931), .ZN(n14095) );
  OR2_X1 U12196 ( .A1(n6575), .A2(n14095), .ZN(n9633) );
  OR2_X1 U12197 ( .A1(n11919), .A2(n9631), .ZN(n9632) );
  NAND4_X1 U12198 ( .A1(n9635), .A2(n9634), .A3(n9633), .A4(n9632), .ZN(n14260) );
  NOR2_X1 U12199 ( .A1(n14883), .A2(n10011), .ZN(n9636) );
  AOI211_X1 U12200 ( .C1(n14217), .C2(n14260), .A(n9637), .B(n9636), .ZN(n9638) );
  OAI211_X1 U12201 ( .C1(n9640), .C2(n14875), .A(n9639), .B(n9638), .ZN(
        P1_U3239) );
  INV_X1 U12202 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10859) );
  XNOR2_X1 U12203 ( .A(n10969), .B(n10859), .ZN(n9643) );
  AOI21_X1 U12204 ( .B1(n10837), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9641), .ZN(
        n9642) );
  NAND2_X1 U12205 ( .A1(n9643), .A2(n9642), .ZN(n10472) );
  OAI21_X1 U12206 ( .B1(n9643), .B2(n9642), .A(n10472), .ZN(n9653) );
  OAI21_X1 U12207 ( .B1(n9645), .B2(n10855), .A(n9644), .ZN(n9647) );
  INV_X1 U12208 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10856) );
  MUX2_X1 U12209 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n10856), .S(n10969), .Z(
        n9646) );
  NAND2_X1 U12210 ( .A1(n9646), .A2(n9647), .ZN(n10478) );
  OAI211_X1 U12211 ( .C1(n9647), .C2(n9646), .A(n14318), .B(n10478), .ZN(n9650) );
  NOR2_X1 U12212 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14112), .ZN(n9648) );
  AOI21_X1 U12213 ( .B1(n14891), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n9648), .ZN(
        n9649) );
  OAI211_X1 U12214 ( .C1(n14320), .C2(n9651), .A(n9650), .B(n9649), .ZN(n9652)
         );
  AOI21_X1 U12215 ( .B1(n14901), .B2(n9653), .A(n9652), .ZN(n9654) );
  INV_X1 U12216 ( .A(n9654), .ZN(P1_U3257) );
  OAI22_X1 U12217 ( .A1(n9671), .A2(n9656), .B1(n9787), .B2(n9655), .ZN(n9658)
         );
  INV_X1 U12218 ( .A(n9671), .ZN(n9666) );
  NAND3_X1 U12219 ( .A1(n9661), .A2(n9660), .A3(n9659), .ZN(n9662) );
  AOI21_X1 U12220 ( .B1(n9787), .B2(n9663), .A(n9662), .ZN(n9664) );
  OAI21_X1 U12221 ( .B1(n9666), .B2(n9665), .A(n9664), .ZN(n9667) );
  NAND2_X1 U12222 ( .A1(n9667), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9670) );
  NAND2_X1 U12223 ( .A1(n9787), .A2(n9668), .ZN(n9669) );
  INV_X1 U12224 ( .A(n12729), .ZN(n12706) );
  NAND2_X1 U12225 ( .A1(n12706), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9826) );
  NAND2_X1 U12226 ( .A1(n9826), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9677) );
  NAND2_X1 U12227 ( .A1(n9671), .A2(n15200), .ZN(n9673) );
  NAND2_X1 U12228 ( .A1(n9786), .A2(n15195), .ZN(n9674) );
  AOI22_X1 U12229 ( .A1(n12737), .A2(n9675), .B1(n12717), .B2(n15173), .ZN(
        n9676) );
  OAI211_X1 U12230 ( .C1(n12930), .C2(n12739), .A(n9677), .B(n9676), .ZN(
        P3_U3172) );
  XNOR2_X1 U12231 ( .A(n11973), .B(n14262), .ZN(n12134) );
  INV_X1 U12232 ( .A(n9678), .ZN(n9679) );
  XOR2_X1 U12233 ( .A(n9922), .B(n12134), .Z(n9740) );
  NAND2_X1 U12234 ( .A1(n14263), .A2(n11966), .ZN(n9682) );
  NAND2_X1 U12235 ( .A1(n9683), .A2(n9682), .ZN(n9685) );
  OR2_X1 U12236 ( .A1(n14263), .A2(n11966), .ZN(n9684) );
  XOR2_X1 U12237 ( .A(n12134), .B(n9940), .Z(n9686) );
  OAI222_X1 U12238 ( .A1(n14637), .A2(n9941), .B1(n14517), .B2(n11965), .C1(
        n14724), .C2(n9686), .ZN(n9737) );
  INV_X1 U12239 ( .A(n9737), .ZN(n9687) );
  MUX2_X1 U12240 ( .A(n9688), .B(n9687), .S(n14544), .Z(n9694) );
  OR2_X1 U12241 ( .A1(n9690), .A2(n11973), .ZN(n10008) );
  INV_X1 U12242 ( .A(n10008), .ZN(n9689) );
  AOI211_X1 U12243 ( .C1(n11973), .C2(n9690), .A(n14924), .B(n9689), .ZN(n9738) );
  OAI22_X1 U12244 ( .A1(n14506), .A2(n7091), .B1(n9691), .B2(n14541), .ZN(
        n9692) );
  AOI21_X1 U12245 ( .B1(n9738), .B2(n14739), .A(n9692), .ZN(n9693) );
  OAI211_X1 U12246 ( .C1(n9740), .C2(n14546), .A(n9694), .B(n9693), .ZN(
        P1_U3288) );
  XNOR2_X1 U12247 ( .A(n13414), .B(n13424), .ZN(n9749) );
  NAND2_X1 U12248 ( .A1(n13555), .A2(n13845), .ZN(n9698) );
  NAND2_X1 U12249 ( .A1(n9747), .A2(n9695), .ZN(n9696) );
  NAND2_X1 U12250 ( .A1(n13554), .A2(n13845), .ZN(n9704) );
  INV_X1 U12251 ( .A(n9749), .ZN(n9700) );
  INV_X1 U12252 ( .A(n9698), .ZN(n9699) );
  NAND2_X1 U12253 ( .A1(n9700), .A2(n9699), .ZN(n9746) );
  NAND2_X1 U12254 ( .A1(n9747), .A2(n9745), .ZN(n9701) );
  INV_X1 U12255 ( .A(n9703), .ZN(n9721) );
  AOI22_X1 U12256 ( .A1(n11505), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n11504), 
        .B2(n9705), .ZN(n9706) );
  NAND2_X1 U12257 ( .A1(n13553), .A2(n13845), .ZN(n9845) );
  NAND2_X1 U12258 ( .A1(n12390), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9714) );
  INV_X1 U12259 ( .A(n9709), .ZN(n9708) );
  NAND2_X1 U12260 ( .A1(n9708), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9859) );
  NAND2_X1 U12261 ( .A1(n9709), .A2(n9867), .ZN(n9710) );
  AND2_X1 U12262 ( .A1(n9859), .A2(n9710), .ZN(n10589) );
  NAND2_X1 U12263 ( .A1(n6638), .A2(n10589), .ZN(n9713) );
  NAND2_X1 U12264 ( .A1(n11618), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9712) );
  NAND2_X1 U12265 ( .A1(n11619), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9711) );
  NAND4_X1 U12266 ( .A1(n9714), .A2(n9713), .A3(n9712), .A4(n9711), .ZN(n13552) );
  NAND2_X1 U12267 ( .A1(n13517), .A2(n13552), .ZN(n9716) );
  NAND2_X1 U12268 ( .A1(n13554), .A2(n13518), .ZN(n9715) );
  AND2_X1 U12269 ( .A1(n9716), .A2(n9715), .ZN(n9767) );
  INV_X1 U12270 ( .A(n13495), .ZN(n13522) );
  NAND2_X1 U12271 ( .A1(n13522), .A2(n9811), .ZN(n9718) );
  OAI211_X1 U12272 ( .C1(n9767), .C2(n13503), .A(n9718), .B(n9717), .ZN(n9719)
         );
  AOI21_X1 U12273 ( .B1(n12259), .B2(n13510), .A(n9719), .ZN(n9724) );
  INV_X1 U12274 ( .A(n13554), .ZN(n9763) );
  OAI22_X1 U12275 ( .A1(n13512), .A2(n9763), .B1(n9721), .B2(n13478), .ZN(
        n9722) );
  NAND3_X1 U12276 ( .A1(n9720), .A2(n6421), .A3(n9722), .ZN(n9723) );
  OAI211_X1 U12277 ( .C1(n9848), .C2(n13478), .A(n9724), .B(n9723), .ZN(
        P2_U3203) );
  INV_X1 U12278 ( .A(n9726), .ZN(n9727) );
  AOI21_X1 U12279 ( .B1(n9728), .B2(n9725), .A(n9727), .ZN(n9736) );
  INV_X1 U12280 ( .A(n9729), .ZN(n9730) );
  OAI22_X1 U12281 ( .A1(n13525), .A2(n12194), .B1(n9730), .B2(n13503), .ZN(
        n9731) );
  AOI21_X1 U12282 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n9837), .A(n9731), .ZN(
        n9735) );
  INV_X1 U12283 ( .A(n13512), .ZN(n13436) );
  INV_X1 U12284 ( .A(n9732), .ZN(n9733) );
  NAND3_X1 U12285 ( .A1(n13436), .A2(n9725), .A3(n9733), .ZN(n9734) );
  OAI211_X1 U12286 ( .C1(n9736), .C2(n13478), .A(n9735), .B(n9734), .ZN(
        P2_U3194) );
  INV_X1 U12287 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9742) );
  AOI211_X1 U12288 ( .C1(n11973), .C2(n14961), .A(n9738), .B(n9737), .ZN(n9739) );
  OAI21_X1 U12289 ( .B1(n14969), .B2(n9740), .A(n9739), .ZN(n9743) );
  NAND2_X1 U12290 ( .A1(n9743), .A2(n14953), .ZN(n9741) );
  OAI21_X1 U12291 ( .B1(n14953), .B2(n9742), .A(n9741), .ZN(P1_U3474) );
  NAND2_X1 U12292 ( .A1(n9743), .A2(n14986), .ZN(n9744) );
  OAI21_X1 U12293 ( .B1(n14986), .B2(n9254), .A(n9744), .ZN(P1_U3533) );
  INV_X1 U12294 ( .A(n9745), .ZN(n9748) );
  NAND2_X1 U12295 ( .A1(n9747), .A2(n9746), .ZN(n13405) );
  AOI21_X1 U12296 ( .B1(n13406), .B2(n9748), .A(n13405), .ZN(n13407) );
  NOR3_X1 U12297 ( .A1(n13512), .A2(n9750), .A3(n9749), .ZN(n9751) );
  AOI21_X1 U12298 ( .B1(n13407), .B2(n13527), .A(n9751), .ZN(n9759) );
  NAND2_X1 U12299 ( .A1(n13521), .A2(n9752), .ZN(n9753) );
  NAND2_X1 U12300 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n15032) );
  OAI211_X1 U12301 ( .C1(n13525), .C2(n9754), .A(n9753), .B(n15032), .ZN(n9756) );
  NOR2_X1 U12302 ( .A1(n9720), .A2(n13478), .ZN(n9755) );
  AOI211_X1 U12303 ( .C1(n13522), .C2(n9996), .A(n9756), .B(n9755), .ZN(n9757)
         );
  OAI21_X1 U12304 ( .B1(n9759), .B2(n9758), .A(n9757), .ZN(P2_U3193) );
  XNOR2_X1 U12305 ( .A(n9907), .B(n12460), .ZN(n9806) );
  AOI21_X1 U12306 ( .B1(n9761), .B2(n12259), .A(n13777), .ZN(n9762) );
  AND2_X1 U12307 ( .A1(n9762), .A2(n9910), .ZN(n9809) );
  OR2_X1 U12308 ( .A1(n12245), .A2(n9763), .ZN(n9764) );
  OAI211_X1 U12309 ( .C1(n9766), .C2(n12460), .A(n9913), .B(n13891), .ZN(n9768) );
  NAND2_X1 U12310 ( .A1(n9768), .A2(n9767), .ZN(n9816) );
  AOI211_X1 U12311 ( .C1(n14012), .C2(n9806), .A(n9809), .B(n9816), .ZN(n9773)
         );
  AOI22_X1 U12312 ( .A1(n13992), .A2(n12259), .B1(n15109), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n9769) );
  OAI21_X1 U12313 ( .B1(n9773), .B2(n15109), .A(n9769), .ZN(P2_U3508) );
  INV_X1 U12314 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9770) );
  NOR2_X1 U12315 ( .A1(n15106), .A2(n9770), .ZN(n9771) );
  AOI21_X1 U12316 ( .B1(n14051), .B2(n12259), .A(n9771), .ZN(n9772) );
  OAI21_X1 U12317 ( .B1(n9773), .B2(n15104), .A(n9772), .ZN(P2_U3457) );
  OAI21_X1 U12318 ( .B1(n9776), .B2(n12773), .A(n9775), .ZN(n9777) );
  XNOR2_X1 U12319 ( .A(n10055), .B(n7722), .ZN(n10056) );
  XNOR2_X1 U12320 ( .A(n10056), .B(n15194), .ZN(n10057) );
  NAND2_X1 U12321 ( .A1(n15173), .A2(n9779), .ZN(n9781) );
  OAI21_X1 U12322 ( .B1(n10055), .B2(n9781), .A(n9784), .ZN(n9821) );
  NAND2_X1 U12323 ( .A1(n12548), .A2(n15188), .ZN(n9783) );
  INV_X1 U12324 ( .A(n9784), .ZN(n9785) );
  XOR2_X1 U12325 ( .A(n10057), .B(n10058), .Z(n9791) );
  NAND2_X1 U12326 ( .A1(n9786), .A2(n15192), .ZN(n12960) );
  AOI22_X1 U12327 ( .A1(n12731), .A2(n15173), .B1(n12717), .B2(n15172), .ZN(
        n9788) );
  OAI21_X1 U12328 ( .B1(n7722), .B2(n12720), .A(n9788), .ZN(n9789) );
  AOI21_X1 U12329 ( .B1(n9826), .B2(P3_REG3_REG_2__SCAN_IN), .A(n9789), .ZN(
        n9790) );
  OAI21_X1 U12330 ( .B1(n9791), .B2(n12739), .A(n9790), .ZN(P3_U3177) );
  INV_X1 U12331 ( .A(n9792), .ZN(n9799) );
  INV_X1 U12332 ( .A(n9793), .ZN(n9796) );
  NAND2_X1 U12333 ( .A1(n13386), .A2(n9794), .ZN(n9795) );
  OAI21_X1 U12334 ( .B1(n13386), .B2(n9796), .A(n9795), .ZN(n9797) );
  INV_X1 U12335 ( .A(n9797), .ZN(n9798) );
  INV_X1 U12336 ( .A(n10287), .ZN(n9801) );
  AOI21_X1 U12337 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n15201), .A(n9801), .ZN(
        n9803) );
  MUX2_X1 U12338 ( .A(n9804), .B(n9803), .S(n15204), .Z(n9805) );
  OAI21_X1 U12339 ( .B1(n12771), .B2(n15165), .A(n9805), .ZN(P3_U3233) );
  INV_X1 U12340 ( .A(n9806), .ZN(n9818) );
  AND2_X1 U12341 ( .A1(n6597), .A2(n9807), .ZN(n9808) );
  NAND2_X1 U12342 ( .A1(n13923), .A2(n9809), .ZN(n9814) );
  NOR2_X2 U12343 ( .A1(n15075), .A2(n9810), .ZN(n13927) );
  NAND2_X1 U12344 ( .A1(n13927), .A2(n12259), .ZN(n9813) );
  AOI22_X1 U12345 ( .A1(n15075), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n9811), .B2(
        n15062), .ZN(n9812) );
  NAND3_X1 U12346 ( .A1(n9814), .A2(n9813), .A3(n9812), .ZN(n9815) );
  AOI21_X1 U12347 ( .B1(n9816), .B2(n13868), .A(n9815), .ZN(n9817) );
  OAI21_X1 U12348 ( .B1(n9818), .B2(n13871), .A(n9817), .ZN(P2_U3256) );
  NOR3_X1 U12349 ( .A1(n15189), .A2(n12548), .A3(n15190), .ZN(n9820) );
  AOI211_X1 U12350 ( .C1(n9822), .C2(n9821), .A(n9820), .B(n9819), .ZN(n9828)
         );
  NOR2_X1 U12351 ( .A1(n12720), .A2(n15187), .ZN(n9825) );
  INV_X1 U12352 ( .A(n15193), .ZN(n9823) );
  OAI22_X1 U12353 ( .A1(n10062), .A2(n12734), .B1(n12719), .B2(n9823), .ZN(
        n9824) );
  AOI211_X1 U12354 ( .C1(n9826), .C2(P3_REG3_REG_1__SCAN_IN), .A(n9825), .B(
        n9824), .ZN(n9827) );
  OAI21_X1 U12355 ( .B1(n9828), .B2(n12739), .A(n9827), .ZN(P3_U3162) );
  INV_X1 U12356 ( .A(n9829), .ZN(n9832) );
  OAI22_X1 U12357 ( .A1(n9830), .A2(P3_U3151), .B1(SI_22_), .B2(n9579), .ZN(
        n9831) );
  AOI21_X1 U12358 ( .B1(n9832), .B2(n13393), .A(n9831), .ZN(P3_U3273) );
  NAND2_X1 U12359 ( .A1(n13436), .A2(n13563), .ZN(n9836) );
  AOI21_X1 U12360 ( .B1(n13777), .B2(n13563), .A(n13478), .ZN(n9833) );
  NOR2_X1 U12361 ( .A1(n9833), .A2(n13510), .ZN(n9835) );
  MUX2_X1 U12362 ( .A(n9836), .B(n9835), .S(n9834), .Z(n9839) );
  NAND2_X1 U12363 ( .A1(n9837), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9838) );
  OAI211_X1 U12364 ( .C1(n13503), .C2(n9840), .A(n9839), .B(n9838), .ZN(
        P2_U3204) );
  AOI22_X1 U12365 ( .A1(n11505), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n11504), 
        .B2(n9841), .ZN(n9842) );
  INV_X1 U12366 ( .A(n9844), .ZN(n9846) );
  NAND2_X1 U12367 ( .A1(n9846), .A2(n9845), .ZN(n9847) );
  AND2_X1 U12368 ( .A1(n13552), .A2(n6649), .ZN(n9849) );
  NAND2_X1 U12369 ( .A1(n11742), .A2(n9849), .ZN(n10206) );
  INV_X1 U12370 ( .A(n11742), .ZN(n9851) );
  INV_X1 U12371 ( .A(n9849), .ZN(n9850) );
  NAND2_X1 U12372 ( .A1(n9851), .A2(n9850), .ZN(n9852) );
  NAND2_X1 U12373 ( .A1(n10206), .A2(n9852), .ZN(n9854) );
  AOI21_X1 U12374 ( .B1(n9853), .B2(n9854), .A(n13478), .ZN(n9857) );
  INV_X1 U12375 ( .A(n9854), .ZN(n9855) );
  NAND2_X1 U12376 ( .A1(n9857), .A2(n11744), .ZN(n9870) );
  INV_X1 U12377 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9858) );
  NAND2_X1 U12378 ( .A1(n9859), .A2(n9858), .ZN(n9860) );
  AND2_X1 U12379 ( .A1(n10214), .A2(n9860), .ZN(n11747) );
  NAND2_X1 U12380 ( .A1(n6638), .A2(n11747), .ZN(n9864) );
  NAND2_X1 U12381 ( .A1(n12390), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9863) );
  NAND2_X1 U12382 ( .A1(n11619), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n9862) );
  NAND2_X1 U12383 ( .A1(n11618), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9861) );
  NAND4_X1 U12384 ( .A1(n9864), .A2(n9863), .A3(n9862), .A4(n9861), .ZN(n13551) );
  NAND2_X1 U12385 ( .A1(n13517), .A2(n13551), .ZN(n9866) );
  NAND2_X1 U12386 ( .A1(n13553), .A2(n13518), .ZN(n9865) );
  AND2_X1 U12387 ( .A1(n9866), .A2(n9865), .ZN(n9915) );
  OAI22_X1 U12388 ( .A1(n13503), .A2(n9915), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9867), .ZN(n9868) );
  AOI21_X1 U12389 ( .B1(n10589), .B2(n13522), .A(n9868), .ZN(n9869) );
  OAI211_X1 U12390 ( .C1(n6950), .C2(n13525), .A(n9870), .B(n9869), .ZN(
        P2_U3189) );
  INV_X1 U12391 ( .A(n11895), .ZN(n9871) );
  NAND2_X1 U12392 ( .A1(n7856), .A2(n9871), .ZN(n10039) );
  NAND2_X1 U12393 ( .A1(n9876), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9874) );
  NAND2_X1 U12394 ( .A1(n7711), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9873) );
  NAND2_X1 U12395 ( .A1(n7852), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9872) );
  INV_X2 U12396 ( .A(P3_U3897), .ZN(n12976) );
  NAND2_X1 U12397 ( .A1(n12976), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n9875) );
  OAI21_X1 U12398 ( .B1(n12755), .B2(n12976), .A(n9875), .ZN(P3_U3521) );
  NAND2_X1 U12399 ( .A1(n9876), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n9879) );
  NAND2_X1 U12400 ( .A1(n10035), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n9878) );
  NAND2_X1 U12401 ( .A1(n7852), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n9877) );
  NAND2_X1 U12402 ( .A1(n12976), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(n9880) );
  OAI21_X1 U12403 ( .B1(n13081), .B2(n12976), .A(n9880), .ZN(P3_U3522) );
  INV_X1 U12404 ( .A(n9888), .ZN(n9883) );
  INV_X1 U12405 ( .A(n9329), .ZN(n9882) );
  INV_X1 U12406 ( .A(n9881), .ZN(n10135) );
  AOI21_X1 U12407 ( .B1(n9883), .B2(n9882), .A(n10135), .ZN(n9895) );
  NAND2_X1 U12408 ( .A1(n13517), .A2(n13557), .ZN(n9885) );
  NAND2_X1 U12409 ( .A1(n13559), .A2(n13518), .ZN(n9884) );
  NAND2_X1 U12410 ( .A1(n9885), .A2(n9884), .ZN(n10303) );
  INV_X1 U12411 ( .A(n10303), .ZN(n9887) );
  NAND2_X1 U12412 ( .A1(n13510), .A2(n15089), .ZN(n9886) );
  NAND2_X1 U12413 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n15001) );
  OAI211_X1 U12414 ( .C1(n9887), .C2(n13503), .A(n9886), .B(n15001), .ZN(n9892) );
  NOR4_X1 U12415 ( .A1(n13512), .A2(n9890), .A3(n9889), .A4(n9888), .ZN(n9891)
         );
  AOI211_X1 U12416 ( .C1(n13522), .C2(n9893), .A(n9892), .B(n9891), .ZN(n9894)
         );
  OAI21_X1 U12417 ( .B1(n9895), .B2(n13478), .A(n9894), .ZN(P2_U3202) );
  INV_X1 U12418 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n13683) );
  NAND2_X1 U12419 ( .A1(n12897), .A2(P3_U3897), .ZN(n9896) );
  OAI21_X1 U12420 ( .B1(P3_U3897), .B2(n13683), .A(n9896), .ZN(P3_U3518) );
  OAI21_X1 U12421 ( .B1(n10210), .B2(P2_REG2_REG_12__SCAN_IN), .A(n9897), .ZN(
        n15055) );
  INV_X1 U12422 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n13725) );
  MUX2_X1 U12423 ( .A(n13725), .B(P2_REG2_REG_13__SCAN_IN), .S(n15051), .Z(
        n15056) );
  NOR2_X1 U12424 ( .A1(n15055), .A2(n15056), .ZN(n15053) );
  XNOR2_X1 U12425 ( .A(n10461), .B(n10460), .ZN(n10462) );
  XNOR2_X1 U12426 ( .A(n10462), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n9905) );
  NOR2_X1 U12427 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11706), .ZN(n9898) );
  AOI21_X1 U12428 ( .B1(n14987), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n9898), .ZN(
        n9899) );
  OAI21_X1 U12429 ( .B1(n10460), .B2(n14993), .A(n9899), .ZN(n9904) );
  OAI21_X1 U12430 ( .B1(n10210), .B2(P2_REG1_REG_12__SCAN_IN), .A(n9900), .ZN(
        n15047) );
  XNOR2_X1 U12431 ( .A(n15051), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n15048) );
  XNOR2_X1 U12432 ( .A(n10648), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n9901) );
  NOR2_X1 U12433 ( .A1(n9902), .A2(n9901), .ZN(n10457) );
  AOI211_X1 U12434 ( .C1(n9902), .C2(n9901), .A(n15046), .B(n10457), .ZN(n9903) );
  AOI211_X1 U12435 ( .C1(n15039), .C2(n9905), .A(n9904), .B(n9903), .ZN(n9906)
         );
  INV_X1 U12436 ( .A(n9906), .ZN(P2_U3228) );
  NAND2_X1 U12437 ( .A1(n9907), .A2(n7197), .ZN(n9909) );
  NAND2_X1 U12438 ( .A1(n12259), .A2(n13553), .ZN(n9908) );
  XNOR2_X1 U12439 ( .A(n12268), .B(n13552), .ZN(n12462) );
  XNOR2_X1 U12440 ( .A(n10238), .B(n12462), .ZN(n10587) );
  AOI21_X1 U12441 ( .B1(n12268), .B2(n9910), .A(n13777), .ZN(n9911) );
  AND2_X1 U12442 ( .A1(n9911), .A2(n10252), .ZN(n10588) );
  INV_X1 U12443 ( .A(n13553), .ZN(n12261) );
  OR2_X1 U12444 ( .A1(n12259), .A2(n12261), .ZN(n9912) );
  OAI211_X1 U12445 ( .C1(n9914), .C2(n12462), .A(n10245), .B(n13891), .ZN(
        n9916) );
  NAND2_X1 U12446 ( .A1(n9916), .A2(n9915), .ZN(n10593) );
  AOI211_X1 U12447 ( .C1(n14012), .C2(n10587), .A(n10588), .B(n10593), .ZN(
        n9921) );
  INV_X1 U12448 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9917) );
  NOR2_X1 U12449 ( .A1(n15106), .A2(n9917), .ZN(n9918) );
  AOI21_X1 U12450 ( .B1(n14051), .B2(n12268), .A(n9918), .ZN(n9919) );
  OAI21_X1 U12451 ( .B1(n9921), .B2(n15104), .A(n9919), .ZN(P2_U3460) );
  AOI22_X1 U12452 ( .A1(n13992), .A2(n12268), .B1(n15109), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n9920) );
  OAI21_X1 U12453 ( .B1(n9921), .B2(n15109), .A(n9920), .ZN(P2_U3509) );
  XNOR2_X1 U12454 ( .A(n14944), .B(n14261), .ZN(n12133) );
  NAND2_X1 U12455 ( .A1(n10005), .A2(n10014), .ZN(n10007) );
  OR2_X1 U12456 ( .A1(n14944), .A2(n14261), .ZN(n9923) );
  NAND2_X1 U12457 ( .A1(n10007), .A2(n9923), .ZN(n9929) );
  OR2_X1 U12458 ( .A1(n9925), .A2(n9924), .ZN(n9928) );
  AOI22_X1 U12459 ( .A1(n12116), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11366), 
        .B2(n9926), .ZN(n9927) );
  XNOR2_X1 U12460 ( .A(n14096), .B(n14260), .ZN(n12136) );
  OAI21_X1 U12461 ( .B1(n9929), .B2(n9944), .A(n10270), .ZN(n9948) );
  INV_X1 U12462 ( .A(n9948), .ZN(n9956) );
  NAND2_X1 U12463 ( .A1(n11459), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9937) );
  INV_X1 U12464 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9930) );
  OR2_X1 U12465 ( .A1(n11921), .A2(n9930), .ZN(n9936) );
  NAND2_X1 U12466 ( .A1(n9931), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10117) );
  OR2_X1 U12467 ( .A1(n9931), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9932) );
  NAND2_X1 U12468 ( .A1(n10117), .A2(n9932), .ZN(n10273) );
  OR2_X1 U12469 ( .A1(n6575), .A2(n10273), .ZN(n9935) );
  OR2_X1 U12470 ( .A1(n11919), .A2(n9933), .ZN(n9934) );
  NAND4_X1 U12471 ( .A1(n9937), .A2(n9936), .A3(n9935), .A4(n9934), .ZN(n14259) );
  OAI22_X1 U12472 ( .A1(n9941), .A2(n14517), .B1(n14869), .B2(n14637), .ZN(
        n9947) );
  AND2_X1 U12473 ( .A1(n9938), .A2(n11973), .ZN(n9939) );
  NAND2_X1 U12474 ( .A1(n14944), .A2(n9941), .ZN(n9943) );
  NAND2_X1 U12475 ( .A1(n9942), .A2(n12136), .ZN(n10276) );
  NAND3_X1 U12476 ( .A1(n10017), .A2(n9944), .A3(n9943), .ZN(n9945) );
  AOI21_X1 U12477 ( .B1(n10276), .B2(n9945), .A(n14724), .ZN(n9946) );
  AOI211_X1 U12478 ( .C1(n14729), .C2(n9948), .A(n9947), .B(n9946), .ZN(n9955)
         );
  MUX2_X1 U12479 ( .A(n9949), .B(n9955), .S(n14544), .Z(n9952) );
  AOI211_X1 U12480 ( .C1(n14096), .C2(n10009), .A(n14924), .B(n10271), .ZN(
        n9953) );
  INV_X1 U12481 ( .A(n14096), .ZN(n10268) );
  OAI22_X1 U12482 ( .A1(n14506), .A2(n10268), .B1(n14095), .B2(n14541), .ZN(
        n9950) );
  AOI21_X1 U12483 ( .B1(n9953), .B2(n14739), .A(n9950), .ZN(n9951) );
  OAI211_X1 U12484 ( .C1(n9956), .C2(n14508), .A(n9952), .B(n9951), .ZN(
        P1_U3286) );
  AOI21_X1 U12485 ( .B1(n14096), .B2(n14961), .A(n9953), .ZN(n9954) );
  OAI211_X1 U12486 ( .C1(n9956), .C2(n14966), .A(n9955), .B(n9954), .ZN(n9958)
         );
  NAND2_X1 U12487 ( .A1(n9958), .A2(n14953), .ZN(n9957) );
  OAI21_X1 U12488 ( .B1(n14953), .B2(n9626), .A(n9957), .ZN(P1_U3480) );
  NAND2_X1 U12489 ( .A1(n9958), .A2(n14986), .ZN(n9959) );
  OAI21_X1 U12490 ( .B1(n14986), .B2(n9631), .A(n9959), .ZN(P1_U3535) );
  AOI22_X1 U12491 ( .A1(n9961), .A2(P3_REG2_REG_5__SCAN_IN), .B1(n9967), .B2(
        n9960), .ZN(n9962) );
  INV_X1 U12492 ( .A(n15127), .ZN(n9977) );
  INV_X1 U12493 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n9963) );
  NAND2_X1 U12494 ( .A1(P3_REG2_REG_7__SCAN_IN), .A2(n9964), .ZN(n10159) );
  OAI21_X1 U12495 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n9964), .A(n10159), .ZN(
        n9993) );
  INV_X1 U12496 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n9965) );
  NOR2_X1 U12497 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9965), .ZN(n10620) );
  AOI21_X1 U12498 ( .B1(n15113), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n10620), .ZN(
        n9974) );
  INV_X1 U12499 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n9970) );
  AOI22_X1 U12500 ( .A1(n9968), .A2(P3_REG1_REG_5__SCAN_IN), .B1(n9967), .B2(
        n9966), .ZN(n15118) );
  MUX2_X1 U12501 ( .A(n9970), .B(P3_REG1_REG_6__SCAN_IN), .S(n15127), .Z(
        n15119) );
  INV_X1 U12502 ( .A(n15117), .ZN(n9969) );
  OAI21_X1 U12503 ( .B1(n9977), .B2(n9970), .A(n9969), .ZN(n10163) );
  OAI21_X1 U12504 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n9971), .A(n10165), .ZN(
        n9972) );
  NAND2_X1 U12505 ( .A1(n9972), .A2(n13023), .ZN(n9973) );
  OAI211_X1 U12506 ( .C1(n15150), .C2(n10164), .A(n9974), .B(n9973), .ZN(n9992) );
  NAND2_X1 U12507 ( .A1(n9976), .A2(n9975), .ZN(n15123) );
  MUX2_X1 U12508 ( .A(n9963), .B(n9970), .S(n13037), .Z(n9978) );
  NAND2_X1 U12509 ( .A1(n9978), .A2(n9977), .ZN(n9981) );
  INV_X1 U12510 ( .A(n9978), .ZN(n9979) );
  NAND2_X1 U12511 ( .A1(n9979), .A2(n15127), .ZN(n9980) );
  NAND2_X1 U12512 ( .A1(n9981), .A2(n9980), .ZN(n15121) );
  AOI21_X1 U12513 ( .B1(n15123), .B2(n15122), .A(n15121), .ZN(n15125) );
  INV_X1 U12514 ( .A(n9981), .ZN(n9989) );
  INV_X1 U12515 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n9983) );
  INV_X1 U12516 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n9982) );
  MUX2_X1 U12517 ( .A(n9983), .B(n9982), .S(n13037), .Z(n9985) );
  NAND2_X1 U12518 ( .A1(n9985), .A2(n9984), .ZN(n10152) );
  INV_X1 U12519 ( .A(n9985), .ZN(n9986) );
  NAND2_X1 U12520 ( .A1(n9986), .A2(n10164), .ZN(n9987) );
  AND2_X1 U12521 ( .A1(n10152), .A2(n9987), .ZN(n9988) );
  OR3_X1 U12522 ( .A1(n15125), .A2(n9989), .A3(n9988), .ZN(n9990) );
  AOI21_X1 U12523 ( .B1(n10153), .B2(n9990), .A(n13078), .ZN(n9991) );
  AOI211_X1 U12524 ( .C1(n15154), .C2(n9993), .A(n9992), .B(n9991), .ZN(n9994)
         );
  INV_X1 U12525 ( .A(n9994), .ZN(P3_U3189) );
  INV_X1 U12526 ( .A(n9995), .ZN(n10002) );
  NAND2_X1 U12527 ( .A1(n13927), .A2(n12245), .ZN(n9998) );
  AOI22_X1 U12528 ( .A1(n15075), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n9996), .B2(
        n15062), .ZN(n9997) );
  NAND2_X1 U12529 ( .A1(n9998), .A2(n9997), .ZN(n10001) );
  NOR2_X1 U12530 ( .A1(n9999), .A2(n13871), .ZN(n10000) );
  AOI211_X1 U12531 ( .C1(n10002), .C2(n13923), .A(n10001), .B(n10000), .ZN(
        n10003) );
  OAI21_X1 U12532 ( .B1(n15075), .B2(n10004), .A(n10003), .ZN(P2_U3257) );
  OR2_X1 U12533 ( .A1(n10005), .A2(n10014), .ZN(n10006) );
  NAND2_X1 U12534 ( .A1(n10007), .A2(n10006), .ZN(n14946) );
  AOI21_X1 U12535 ( .B1(n10008), .B2(n14944), .A(n14924), .ZN(n10010) );
  NAND2_X1 U12536 ( .A1(n10010), .A2(n10009), .ZN(n14947) );
  INV_X1 U12537 ( .A(n10011), .ZN(n10012) );
  AOI22_X1 U12538 ( .A1(n14733), .A2(n14944), .B1(n14732), .B2(n10012), .ZN(
        n10013) );
  OAI21_X1 U12539 ( .B1(n14486), .B2(n14947), .A(n10013), .ZN(n10025) );
  NAND2_X1 U12540 ( .A1(n14946), .A2(n14729), .ZN(n10023) );
  NAND2_X1 U12541 ( .A1(n10015), .A2(n10014), .ZN(n10016) );
  NAND2_X1 U12542 ( .A1(n10017), .A2(n10016), .ZN(n10021) );
  NAND2_X1 U12543 ( .A1(n14262), .A2(n14394), .ZN(n10019) );
  NAND2_X1 U12544 ( .A1(n14260), .A2(n14921), .ZN(n10018) );
  NAND2_X1 U12545 ( .A1(n10019), .A2(n10018), .ZN(n10020) );
  AOI21_X1 U12546 ( .B1(n10021), .B2(n14832), .A(n10020), .ZN(n10022) );
  NAND2_X1 U12547 ( .A1(n10023), .A2(n10022), .ZN(n14951) );
  MUX2_X1 U12548 ( .A(n14951), .B(P1_REG2_REG_6__SCAN_IN), .S(n14743), .Z(
        n10024) );
  AOI211_X1 U12549 ( .C1(n14740), .C2(n14946), .A(n10025), .B(n10024), .ZN(
        n10026) );
  INV_X1 U12550 ( .A(n10026), .ZN(P1_U3287) );
  AOI22_X1 U12551 ( .A1(n13927), .A2(n12227), .B1(n15062), .B2(n10139), .ZN(
        n10027) );
  OAI21_X1 U12552 ( .B1(n13866), .B2(n10028), .A(n10027), .ZN(n10029) );
  AOI21_X1 U12553 ( .B1(n15072), .B2(n10030), .A(n10029), .ZN(n10034) );
  MUX2_X1 U12554 ( .A(n10032), .B(n10031), .S(n15075), .Z(n10033) );
  NAND2_X1 U12555 ( .A1(n10034), .A2(n10033), .ZN(P2_U3260) );
  INV_X1 U12556 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n13673) );
  NAND2_X1 U12557 ( .A1(n10035), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n10038) );
  NAND2_X1 U12558 ( .A1(n7974), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n10037) );
  NAND2_X1 U12559 ( .A1(n7852), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n10036) );
  INV_X1 U12560 ( .A(n13089), .ZN(n10040) );
  NAND2_X1 U12561 ( .A1(n10040), .A2(P3_U3897), .ZN(n10041) );
  OAI21_X1 U12562 ( .B1(P3_U3897), .B2(n13673), .A(n10041), .ZN(P3_U3520) );
  OR2_X1 U12563 ( .A1(n15200), .A2(n10042), .ZN(n15183) );
  NAND2_X1 U12564 ( .A1(n15177), .A2(n15183), .ZN(n14779) );
  OAI21_X1 U12565 ( .B1(n10044), .B2(n12929), .A(n10043), .ZN(n10045) );
  INV_X1 U12566 ( .A(n10045), .ZN(n10068) );
  OAI211_X1 U12567 ( .C1(n10048), .C2(n10047), .A(n10046), .B(n14762), .ZN(
        n10050) );
  AOI22_X1 U12568 ( .A1(n15192), .A2(n15194), .B1(n12975), .B2(n15195), .ZN(
        n10049) );
  AND2_X1 U12569 ( .A1(n10050), .A2(n10049), .ZN(n10067) );
  MUX2_X1 U12570 ( .A(n10067), .B(n10051), .S(n15206), .Z(n10054) );
  INV_X1 U12571 ( .A(n15165), .ZN(n11101) );
  AOI22_X1 U12572 ( .A1(n11101), .A2(n10052), .B1(n15201), .B2(n7724), .ZN(
        n10053) );
  OAI211_X1 U12573 ( .C1(n13207), .C2(n10068), .A(n10054), .B(n10053), .ZN(
        P3_U3230) );
  XNOR2_X1 U12574 ( .A(n10055), .B(n10495), .ZN(n10089) );
  XNOR2_X1 U12575 ( .A(n10089), .B(n15172), .ZN(n10060) );
  INV_X1 U12577 ( .A(n10061), .ZN(n10066) );
  OAI22_X1 U12578 ( .A1(n12720), .A2(n10495), .B1(n10062), .B2(n12719), .ZN(
        n10063) );
  AOI211_X1 U12579 ( .C1(n12717), .C2(n12975), .A(n10064), .B(n10063), .ZN(
        n10065) );
  OAI211_X1 U12580 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12706), .A(n10066), .B(
        n10065), .ZN(P3_U3158) );
  OAI21_X1 U12581 ( .B1(n14790), .B2(n10068), .A(n10067), .ZN(n10497) );
  INV_X1 U12582 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n10069) );
  OAI22_X1 U12583 ( .A1(n10495), .A2(n13384), .B1(n15232), .B2(n10069), .ZN(
        n10070) );
  AOI21_X1 U12584 ( .B1(n10497), .B2(n15232), .A(n10070), .ZN(n10071) );
  INV_X1 U12585 ( .A(n10071), .ZN(P3_U3399) );
  NAND2_X1 U12586 ( .A1(n10072), .A2(n13393), .ZN(n10073) );
  OAI211_X1 U12587 ( .C1(n10074), .C2(n9579), .A(n10073), .B(n12959), .ZN(
        P3_U3272) );
  NAND2_X1 U12588 ( .A1(n10075), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10076) );
  XNOR2_X1 U12589 ( .A(n10076), .B(P2_IR_REG_18__SCAN_IN), .ZN(n11225) );
  INV_X1 U12590 ( .A(n11225), .ZN(n11261) );
  INV_X1 U12591 ( .A(n10079), .ZN(n10081) );
  NAND2_X1 U12592 ( .A1(n10081), .A2(n10080), .ZN(n10082) );
  XNOR2_X1 U12593 ( .A(n10194), .B(SI_18_), .ZN(n10193) );
  MUX2_X1 U12594 ( .A(n10087), .B(n10083), .S(n11907), .Z(n10180) );
  XNOR2_X1 U12595 ( .A(n10193), .B(n10180), .ZN(n11357) );
  INV_X1 U12596 ( .A(n11357), .ZN(n10086) );
  OAI222_X1 U12597 ( .A1(P2_U3088), .A2(n11261), .B1(n14086), .B2(n10083), 
        .C1(n14088), .C2(n10086), .ZN(P2_U3309) );
  OAI21_X1 U12598 ( .B1(n10084), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10085) );
  XNOR2_X1 U12599 ( .A(n10085), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14314) );
  INV_X1 U12600 ( .A(n14314), .ZN(n14307) );
  OAI222_X1 U12601 ( .A1(n14307), .A2(P1_U3086), .B1(n14689), .B2(n10087), 
        .C1(n14694), .C2(n10086), .ZN(P1_U3337) );
  INV_X1 U12602 ( .A(n10088), .ZN(n10437) );
  INV_X4 U12603 ( .A(n12548), .ZN(n12614) );
  XNOR2_X1 U12604 ( .A(n10055), .B(n12787), .ZN(n10260) );
  OAI21_X1 U12605 ( .B1(n10091), .B2(n10090), .A(n10262), .ZN(n10092) );
  NAND2_X1 U12606 ( .A1(n10092), .A2(n12673), .ZN(n10097) );
  OAI22_X1 U12607 ( .A1(n12720), .A2(n12787), .B1(n10093), .B2(n12719), .ZN(
        n10094) );
  AOI211_X1 U12608 ( .C1(n12717), .C2(n12974), .A(n10095), .B(n10094), .ZN(
        n10096) );
  OAI211_X1 U12609 ( .C1(n10437), .C2(n12706), .A(n10097), .B(n10096), .ZN(
        P3_U3170) );
  OR2_X1 U12610 ( .A1(n10098), .A2(n9924), .ZN(n10101) );
  AOI22_X1 U12611 ( .A1(n12116), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11366), 
        .B2(n10099), .ZN(n10100) );
  NAND2_X1 U12612 ( .A1(n10101), .A2(n10100), .ZN(n14956) );
  AOI22_X1 U12613 ( .A1(n14956), .A2(n6423), .B1(n11874), .B2(n14259), .ZN(
        n11005) );
  NAND2_X1 U12614 ( .A1(n14956), .A2(n11870), .ZN(n10103) );
  NAND2_X1 U12615 ( .A1(n14259), .A2(n11825), .ZN(n10102) );
  NAND2_X1 U12616 ( .A1(n10103), .A2(n10102), .ZN(n10104) );
  XNOR2_X1 U12617 ( .A(n10104), .B(n11881), .ZN(n11002) );
  XOR2_X1 U12618 ( .A(n11005), .B(n11002), .Z(n10115) );
  INV_X1 U12619 ( .A(n14260), .ZN(n10274) );
  NOR2_X1 U12620 ( .A1(n10274), .A2(n11879), .ZN(n10105) );
  AOI21_X1 U12621 ( .B1(n14096), .B2(n6423), .A(n10105), .ZN(n10113) );
  NAND2_X1 U12622 ( .A1(n14096), .A2(n11870), .ZN(n10107) );
  NAND2_X1 U12623 ( .A1(n14260), .A2(n11825), .ZN(n10106) );
  NAND2_X1 U12624 ( .A1(n10107), .A2(n10106), .ZN(n10108) );
  XNOR2_X1 U12625 ( .A(n10108), .B(n11881), .ZN(n10111) );
  INV_X1 U12626 ( .A(n10111), .ZN(n10112) );
  XNOR2_X1 U12627 ( .A(n10111), .B(n10113), .ZN(n14093) );
  OAI21_X1 U12628 ( .B1(n10113), .B2(n10112), .A(n14092), .ZN(n10114) );
  AOI21_X1 U12629 ( .B1(n10115), .B2(n10114), .A(n11003), .ZN(n10129) );
  NAND2_X1 U12630 ( .A1(n11381), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10123) );
  NAND2_X1 U12631 ( .A1(n10117), .A2(n10116), .ZN(n10118) );
  NAND2_X1 U12632 ( .A1(n10384), .A2(n10118), .ZN(n14882) );
  OR2_X1 U12633 ( .A1(n6575), .A2(n14882), .ZN(n10122) );
  OR2_X1 U12634 ( .A1(n11919), .A2(n10119), .ZN(n10121) );
  OR2_X1 U12635 ( .A1(n9229), .A2(n10398), .ZN(n10120) );
  NAND4_X1 U12636 ( .A1(n10123), .A2(n10122), .A3(n10121), .A4(n10120), .ZN(
        n14258) );
  INV_X1 U12637 ( .A(n14258), .ZN(n14807) );
  OAI22_X1 U12638 ( .A1(n14871), .A2(n14807), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13634), .ZN(n10124) );
  INV_X1 U12639 ( .A(n10124), .ZN(n10126) );
  NAND2_X1 U12640 ( .A1(n14115), .A2(n14260), .ZN(n10125) );
  OAI211_X1 U12641 ( .C1(n14883), .C2(n10273), .A(n10126), .B(n10125), .ZN(
        n10127) );
  AOI21_X1 U12642 ( .B1(n14879), .B2(n14956), .A(n10127), .ZN(n10128) );
  OAI21_X1 U12643 ( .B1(n10129), .B2(n14875), .A(n10128), .ZN(P1_U3221) );
  INV_X1 U12644 ( .A(n10130), .ZN(n10132) );
  NAND2_X1 U12645 ( .A1(n13510), .A2(n12227), .ZN(n10131) );
  NAND2_X1 U12646 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n15020) );
  OAI211_X1 U12647 ( .C1(n10132), .C2(n13503), .A(n10131), .B(n15020), .ZN(
        n10138) );
  AOI22_X1 U12648 ( .A1(n13436), .A2(n13558), .B1(n13527), .B2(n10133), .ZN(
        n10136) );
  NOR3_X1 U12649 ( .A1(n10136), .A2(n10135), .A3(n10134), .ZN(n10137) );
  AOI211_X1 U12650 ( .C1(n13522), .C2(n10139), .A(n10138), .B(n10137), .ZN(
        n10140) );
  OAI21_X1 U12651 ( .B1(n10141), .B2(n13478), .A(n10140), .ZN(P2_U3199) );
  OAI21_X1 U12652 ( .B1(n10143), .B2(n12937), .A(n10142), .ZN(n10441) );
  OAI211_X1 U12653 ( .C1(n10146), .C2(n10145), .A(n10144), .B(n14762), .ZN(
        n10148) );
  AOI22_X1 U12654 ( .A1(n15195), .A2(n12974), .B1(n15172), .B2(n15192), .ZN(
        n10147) );
  NAND2_X1 U12655 ( .A1(n10148), .A2(n10147), .ZN(n10438) );
  AOI21_X1 U12656 ( .B1(n14798), .B2(n10441), .A(n10438), .ZN(n10493) );
  INV_X1 U12657 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n10149) );
  OAI22_X1 U12658 ( .A1(n12787), .A2(n13384), .B1(n15232), .B2(n10149), .ZN(
        n10150) );
  INV_X1 U12659 ( .A(n10150), .ZN(n10151) );
  OAI21_X1 U12660 ( .B1(n10493), .B2(n15234), .A(n10151), .ZN(P3_U3402) );
  MUX2_X1 U12661 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13037), .Z(n10154) );
  NAND2_X1 U12662 ( .A1(n10153), .A2(n10152), .ZN(n15145) );
  XOR2_X1 U12663 ( .A(n15149), .B(n10154), .Z(n15144) );
  NAND2_X1 U12664 ( .A1(n15145), .A2(n15144), .ZN(n15143) );
  MUX2_X1 U12665 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n13037), .Z(n10155) );
  NOR2_X1 U12666 ( .A1(n10155), .A2(n10343), .ZN(n10333) );
  INV_X1 U12667 ( .A(n10333), .ZN(n10156) );
  NAND2_X1 U12668 ( .A1(n10155), .A2(n10343), .ZN(n10334) );
  NAND2_X1 U12669 ( .A1(n10156), .A2(n10334), .ZN(n10157) );
  XNOR2_X1 U12670 ( .A(n10335), .B(n10157), .ZN(n10176) );
  NAND2_X1 U12671 ( .A1(n10164), .A2(n10158), .ZN(n10160) );
  INV_X1 U12672 ( .A(n15149), .ZN(n10168) );
  INV_X1 U12673 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10161) );
  NAND2_X1 U12674 ( .A1(P3_REG2_REG_9__SCAN_IN), .A2(n10162), .ZN(n10337) );
  OAI21_X1 U12675 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n10162), .A(n10337), .ZN(
        n10174) );
  INV_X1 U12676 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15238) );
  NAND2_X1 U12677 ( .A1(n10164), .A2(n10163), .ZN(n10166) );
  NAND2_X1 U12678 ( .A1(n10166), .A2(n10165), .ZN(n15137) );
  MUX2_X1 U12679 ( .A(n15238), .B(P3_REG1_REG_8__SCAN_IN), .S(n15149), .Z(
        n15138) );
  INV_X1 U12680 ( .A(n15138), .ZN(n10167) );
  NAND2_X1 U12681 ( .A1(n15137), .A2(n10167), .ZN(n15141) );
  OAI21_X1 U12682 ( .B1(n10168), .B2(n15238), .A(n15141), .ZN(n10342) );
  OAI21_X1 U12683 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n10169), .A(n10344), .ZN(
        n10170) );
  NAND2_X1 U12684 ( .A1(n10170), .A2(n13023), .ZN(n10172) );
  AND2_X1 U12685 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n10962) );
  AOI21_X1 U12686 ( .B1(n15113), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n10962), .ZN(
        n10171) );
  OAI211_X1 U12687 ( .C1(n15150), .C2(n10343), .A(n10172), .B(n10171), .ZN(
        n10173) );
  AOI21_X1 U12688 ( .B1(n10174), .B2(n15154), .A(n10173), .ZN(n10175) );
  OAI21_X1 U12689 ( .B1(n10176), .B2(n13078), .A(n10175), .ZN(P3_U3191) );
  INV_X1 U12690 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10192) );
  NAND2_X1 U12691 ( .A1(n10199), .A2(SI_19_), .ZN(n10182) );
  OAI21_X1 U12692 ( .B1(n10177), .B2(n10180), .A(n10182), .ZN(n10178) );
  INV_X1 U12693 ( .A(n10178), .ZN(n10179) );
  INV_X1 U12694 ( .A(n10180), .ZN(n10196) );
  NOR2_X1 U12695 ( .A1(n10196), .A2(SI_18_), .ZN(n10183) );
  INV_X1 U12696 ( .A(n10199), .ZN(n10181) );
  AOI22_X1 U12697 ( .A1(n10183), .A2(n10182), .B1(n10198), .B2(n10181), .ZN(
        n10184) );
  INV_X1 U12698 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11512) );
  MUX2_X1 U12699 ( .A(n10192), .B(n11512), .S(n11907), .Z(n10189) );
  NAND2_X1 U12700 ( .A1(n10190), .A2(n10189), .ZN(n10191) );
  INV_X1 U12701 ( .A(n11511), .ZN(n11474) );
  OAI222_X1 U12702 ( .A1(P1_U3086), .A2(n6699), .B1(n14689), .B2(n10192), .C1(
        n14694), .C2(n11474), .ZN(P1_U3335) );
  INV_X1 U12703 ( .A(n10193), .ZN(n10197) );
  INV_X1 U12704 ( .A(n10194), .ZN(n10195) );
  XNOR2_X1 U12705 ( .A(n10199), .B(n10198), .ZN(n10200) );
  XNOR2_X1 U12706 ( .A(n10201), .B(n10200), .ZN(n11503) );
  INV_X1 U12707 ( .A(n11503), .ZN(n10258) );
  OAI222_X1 U12708 ( .A1(n14088), .A2(n10258), .B1(n14086), .B2(n10202), .C1(
        P2_U3088), .C2(n13574), .ZN(P2_U3308) );
  NAND2_X1 U12709 ( .A1(n10532), .A2(n12393), .ZN(n10205) );
  AOI22_X1 U12710 ( .A1(n11505), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n11504), 
        .B2(n10203), .ZN(n10204) );
  NAND2_X1 U12711 ( .A1(n13551), .A2(n13845), .ZN(n10208) );
  INV_X1 U12712 ( .A(n10230), .ZN(n10209) );
  AOI22_X1 U12713 ( .A1(n11505), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n11504), 
        .B2(n10210), .ZN(n10211) );
  INV_X1 U12714 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n13616) );
  NAND2_X1 U12715 ( .A1(n10214), .A2(n13616), .ZN(n10215) );
  AND2_X1 U12716 ( .A1(n10220), .A2(n10215), .ZN(n10362) );
  NAND2_X1 U12717 ( .A1(n6638), .A2(n10362), .ZN(n10219) );
  NAND2_X1 U12718 ( .A1(n12390), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10218) );
  NAND2_X1 U12719 ( .A1(n11618), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n10217) );
  NAND2_X1 U12720 ( .A1(n11619), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n10216) );
  NAND4_X1 U12721 ( .A1(n10219), .A2(n10218), .A3(n10217), .A4(n10216), .ZN(
        n13550) );
  NAND2_X1 U12722 ( .A1(n13550), .A2(n13845), .ZN(n10407) );
  NAND2_X1 U12723 ( .A1(n10220), .A2(n10426), .ZN(n10221) );
  AND2_X1 U12724 ( .A1(n10418), .A2(n10221), .ZN(n10563) );
  NAND2_X1 U12725 ( .A1(n6638), .A2(n10563), .ZN(n10225) );
  NAND2_X1 U12726 ( .A1(n12390), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10224) );
  NAND2_X1 U12727 ( .A1(n11619), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n10223) );
  NAND2_X1 U12728 ( .A1(n11618), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10222) );
  NAND4_X1 U12729 ( .A1(n10225), .A2(n10224), .A3(n10223), .A4(n10222), .ZN(
        n13549) );
  NAND2_X1 U12730 ( .A1(n13517), .A2(n13549), .ZN(n10227) );
  NAND2_X1 U12731 ( .A1(n13551), .A2(n13518), .ZN(n10226) );
  AND2_X1 U12732 ( .A1(n10227), .A2(n10226), .ZN(n10360) );
  NAND2_X1 U12733 ( .A1(n13522), .A2(n10362), .ZN(n10229) );
  OAI211_X1 U12734 ( .C1(n10360), .C2(n13503), .A(n10229), .B(n10228), .ZN(
        n10235) );
  INV_X1 U12735 ( .A(n11755), .ZN(n10233) );
  AOI22_X1 U12736 ( .A1(n10230), .A2(n13527), .B1(n13436), .B2(n13551), .ZN(
        n10231) );
  NOR3_X1 U12737 ( .A1(n10233), .A2(n10232), .A3(n10231), .ZN(n10234) );
  AOI211_X1 U12738 ( .C1(n6604), .C2(n13510), .A(n10235), .B(n10234), .ZN(
        n10236) );
  OAI21_X1 U12739 ( .B1(n10410), .B2(n13478), .A(n10236), .ZN(P2_U3196) );
  INV_X1 U12740 ( .A(n12462), .ZN(n10237) );
  NAND2_X1 U12741 ( .A1(n10238), .A2(n10237), .ZN(n10240) );
  NAND2_X1 U12742 ( .A1(n12268), .A2(n13552), .ZN(n10239) );
  INV_X1 U12743 ( .A(n13551), .ZN(n10241) );
  NAND2_X1 U12744 ( .A1(n6651), .A2(n10241), .ZN(n10358) );
  OR2_X1 U12745 ( .A1(n6651), .A2(n10241), .ZN(n10242) );
  NAND2_X1 U12746 ( .A1(n10358), .A2(n10242), .ZN(n12464) );
  XNOR2_X1 U12747 ( .A(n10369), .B(n12464), .ZN(n10332) );
  INV_X1 U12748 ( .A(n13552), .ZN(n10243) );
  OR2_X1 U12749 ( .A1(n12268), .A2(n10243), .ZN(n10244) );
  NAND2_X1 U12750 ( .A1(n10245), .A2(n10244), .ZN(n10246) );
  INV_X1 U12751 ( .A(n10246), .ZN(n10248) );
  INV_X1 U12752 ( .A(n12464), .ZN(n10247) );
  OR2_X2 U12753 ( .A1(n10246), .A2(n12464), .ZN(n10359) );
  OAI21_X1 U12754 ( .B1(n10248), .B2(n10247), .A(n10359), .ZN(n10251) );
  NAND2_X1 U12755 ( .A1(n13517), .A2(n13550), .ZN(n10250) );
  NAND2_X1 U12756 ( .A1(n13552), .A2(n13518), .ZN(n10249) );
  NAND2_X1 U12757 ( .A1(n10250), .A2(n10249), .ZN(n11746) );
  AOI21_X1 U12758 ( .B1(n10251), .B2(n13891), .A(n11746), .ZN(n10327) );
  AOI211_X1 U12759 ( .C1(n6651), .C2(n10252), .A(n6649), .B(n10363), .ZN(
        n10330) );
  AOI21_X1 U12760 ( .B1(n15098), .B2(n6651), .A(n10330), .ZN(n10253) );
  OAI211_X1 U12761 ( .C1(n15093), .C2(n10332), .A(n10327), .B(n10253), .ZN(
        n10255) );
  NAND2_X1 U12762 ( .A1(n10255), .A2(n15112), .ZN(n10254) );
  OAI21_X1 U12763 ( .B1(n15112), .B2(n8891), .A(n10254), .ZN(P2_U3510) );
  INV_X1 U12764 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10257) );
  NAND2_X1 U12765 ( .A1(n10255), .A2(n15106), .ZN(n10256) );
  OAI21_X1 U12766 ( .B1(n15106), .B2(n10257), .A(n10256), .ZN(P2_U3463) );
  OAI222_X1 U12767 ( .A1(P1_U3086), .A2(n14540), .B1(n14689), .B2(n10259), 
        .C1(n14694), .C2(n10258), .ZN(P1_U3336) );
  NAND2_X1 U12768 ( .A1(n10262), .A2(n10261), .ZN(n10611) );
  XNOR2_X1 U12769 ( .A(n12614), .B(n10583), .ZN(n10612) );
  XOR2_X1 U12770 ( .A(n12974), .B(n10612), .Z(n10610) );
  XOR2_X1 U12771 ( .A(n10611), .B(n10610), .Z(n10267) );
  OAI22_X1 U12772 ( .A1(n12720), .A2(n10583), .B1(n6635), .B2(n12719), .ZN(
        n10263) );
  AOI211_X1 U12773 ( .C1(n12717), .C2(n12973), .A(n10264), .B(n10263), .ZN(
        n10266) );
  NAND2_X1 U12774 ( .A1(n12729), .A2(n10584), .ZN(n10265) );
  OAI211_X1 U12775 ( .C1(n10267), .C2(n12739), .A(n10266), .B(n10265), .ZN(
        P3_U3167) );
  XNOR2_X1 U12776 ( .A(n14956), .B(n14869), .ZN(n12138) );
  NAND2_X1 U12777 ( .A1(n10268), .A2(n10274), .ZN(n10269) );
  XOR2_X1 U12778 ( .A(n10376), .B(n12138), .Z(n14958) );
  NAND2_X1 U12779 ( .A1(n10271), .A2(n10375), .ZN(n10399) );
  OR2_X1 U12780 ( .A1(n10271), .A2(n10375), .ZN(n10272) );
  AND3_X1 U12781 ( .A1(n10399), .A2(n14736), .A3(n10272), .ZN(n14955) );
  OAI22_X1 U12782 ( .A1(n14506), .A2(n10375), .B1(n14541), .B2(n10273), .ZN(
        n10284) );
  NAND2_X1 U12783 ( .A1(n14096), .A2(n10274), .ZN(n10275) );
  NAND2_X1 U12784 ( .A1(n10276), .A2(n10275), .ZN(n10279) );
  INV_X1 U12785 ( .A(n10279), .ZN(n10278) );
  NAND2_X1 U12786 ( .A1(n10278), .A2(n10277), .ZN(n10392) );
  NAND2_X1 U12787 ( .A1(n10279), .A2(n12138), .ZN(n10280) );
  NAND3_X1 U12788 ( .A1(n10392), .A2(n14832), .A3(n10280), .ZN(n10282) );
  AOI22_X1 U12789 ( .A1(n14394), .A2(n14260), .B1(n14258), .B2(n14921), .ZN(
        n10281) );
  NAND2_X1 U12790 ( .A1(n10282), .A2(n10281), .ZN(n14954) );
  MUX2_X1 U12791 ( .A(n14954), .B(P1_REG2_REG_8__SCAN_IN), .S(n14743), .Z(
        n10283) );
  AOI211_X1 U12792 ( .C1(n14955), .C2(n14739), .A(n10284), .B(n10283), .ZN(
        n10285) );
  OAI21_X1 U12793 ( .B1(n14546), .B2(n14958), .A(n10285), .ZN(P1_U3285) );
  MUX2_X1 U12794 ( .A(n10287), .B(n10286), .S(n15241), .Z(n10288) );
  OAI21_X1 U12795 ( .B1(n12771), .B2(n13334), .A(n10288), .ZN(P3_U3459) );
  OAI21_X1 U12796 ( .B1(n10290), .B2(n12451), .A(n10289), .ZN(n10291) );
  INV_X1 U12797 ( .A(n10291), .ZN(n15092) );
  INV_X1 U12798 ( .A(n10292), .ZN(n10295) );
  INV_X1 U12799 ( .A(n10293), .ZN(n10294) );
  AOI211_X1 U12800 ( .C1(n15089), .C2(n10295), .A(n6649), .B(n10294), .ZN(
        n15088) );
  OAI22_X1 U12801 ( .A1(n15069), .A2(n10297), .B1(n10296), .B2(n13825), .ZN(
        n10298) );
  AOI21_X1 U12802 ( .B1(n15064), .B2(n15088), .A(n10298), .ZN(n10307) );
  NAND3_X1 U12803 ( .A1(n10300), .A2(n12451), .A3(n10299), .ZN(n10301) );
  AOI21_X1 U12804 ( .B1(n10302), .B2(n10301), .A(n13875), .ZN(n10304) );
  NOR2_X1 U12805 ( .A1(n10304), .A2(n10303), .ZN(n15090) );
  MUX2_X1 U12806 ( .A(n15090), .B(n10305), .S(n15075), .Z(n10306) );
  OAI211_X1 U12807 ( .C1(n15092), .C2(n13871), .A(n10307), .B(n10306), .ZN(
        P2_U3261) );
  OAI21_X1 U12808 ( .B1(n10309), .B2(n7209), .A(n10308), .ZN(n10310) );
  INV_X1 U12809 ( .A(n10310), .ZN(n15102) );
  OAI21_X1 U12810 ( .B1(n10312), .B2(n12456), .A(n10311), .ZN(n10316) );
  NOR2_X1 U12811 ( .A1(n15102), .A2(n6597), .ZN(n10314) );
  AOI211_X1 U12812 ( .C1(n13891), .C2(n10316), .A(n10315), .B(n10314), .ZN(
        n15100) );
  MUX2_X1 U12813 ( .A(n10317), .B(n15100), .S(n13868), .Z(n10324) );
  AOI211_X1 U12814 ( .C1(n15097), .C2(n10319), .A(n6649), .B(n10318), .ZN(
        n15096) );
  INV_X1 U12815 ( .A(n15097), .ZN(n10321) );
  OAI22_X1 U12816 ( .A1(n15069), .A2(n10321), .B1(n10320), .B2(n13825), .ZN(
        n10322) );
  AOI21_X1 U12817 ( .B1(n15064), .B2(n15096), .A(n10322), .ZN(n10323) );
  OAI211_X1 U12818 ( .C1(n15102), .C2(n10325), .A(n10324), .B(n10323), .ZN(
        P2_U3259) );
  INV_X1 U12819 ( .A(n6651), .ZN(n11750) );
  AOI22_X1 U12820 ( .A1(n15075), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11747), 
        .B2(n15062), .ZN(n10326) );
  OAI21_X1 U12821 ( .B1(n11750), .B2(n15069), .A(n10326), .ZN(n10329) );
  NOR2_X1 U12822 ( .A1(n10327), .A2(n15075), .ZN(n10328) );
  AOI211_X1 U12823 ( .C1(n10330), .C2(n15064), .A(n10329), .B(n10328), .ZN(
        n10331) );
  OAI21_X1 U12824 ( .B1(n13871), .B2(n10332), .A(n10331), .ZN(P2_U3254) );
  MUX2_X1 U12825 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13037), .Z(n10502) );
  XOR2_X1 U12826 ( .A(n10346), .B(n10502), .Z(n10503) );
  AOI21_X1 U12827 ( .B1(n10335), .B2(n10334), .A(n10333), .ZN(n10504) );
  XOR2_X1 U12828 ( .A(n10503), .B(n10504), .Z(n10357) );
  NAND2_X1 U12829 ( .A1(n10343), .A2(n10336), .ZN(n10338) );
  NAND2_X1 U12830 ( .A1(n10338), .A2(n10337), .ZN(n10341) );
  INV_X1 U12831 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10339) );
  MUX2_X1 U12832 ( .A(n10339), .B(P3_REG2_REG_10__SCAN_IN), .S(n10346), .Z(
        n10340) );
  NAND2_X1 U12833 ( .A1(n10340), .A2(n10341), .ZN(n10505) );
  OAI21_X1 U12834 ( .B1(n10341), .B2(n10340), .A(n10505), .ZN(n10355) );
  NAND2_X1 U12835 ( .A1(n10343), .A2(n10342), .ZN(n10345) );
  NAND2_X1 U12836 ( .A1(n10345), .A2(n10344), .ZN(n10349) );
  INV_X1 U12837 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n10347) );
  MUX2_X1 U12838 ( .A(n10347), .B(P3_REG1_REG_10__SCAN_IN), .S(n10346), .Z(
        n10348) );
  NAND2_X1 U12839 ( .A1(n10348), .A2(n10349), .ZN(n10509) );
  OAI21_X1 U12840 ( .B1(n10349), .B2(n10348), .A(n10509), .ZN(n10350) );
  NAND2_X1 U12841 ( .A1(n10350), .A2(n13023), .ZN(n10353) );
  NAND2_X1 U12842 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n12589)
         );
  INV_X1 U12843 ( .A(n12589), .ZN(n10351) );
  AOI21_X1 U12844 ( .B1(n15113), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n10351), 
        .ZN(n10352) );
  OAI211_X1 U12845 ( .C1(n15150), .C2(n10508), .A(n10353), .B(n10352), .ZN(
        n10354) );
  AOI21_X1 U12846 ( .B1(n10355), .B2(n15154), .A(n10354), .ZN(n10356) );
  OAI21_X1 U12847 ( .B1(n10357), .B2(n13078), .A(n10356), .ZN(P3_U3192) );
  XNOR2_X1 U12848 ( .A(n12281), .B(n13550), .ZN(n12466) );
  INV_X1 U12849 ( .A(n12466), .ZN(n10566) );
  OAI211_X1 U12850 ( .C1(n6547), .C2(n12466), .A(n13891), .B(n10559), .ZN(
        n10361) );
  NAND2_X1 U12851 ( .A1(n10361), .A2(n10360), .ZN(n10431) );
  AOI21_X1 U12852 ( .B1(n10362), .B2(n15062), .A(n10431), .ZN(n10374) );
  INV_X1 U12853 ( .A(n10363), .ZN(n10365) );
  INV_X1 U12854 ( .A(n6604), .ZN(n10367) );
  INV_X1 U12855 ( .A(n10562), .ZN(n10364) );
  AOI211_X1 U12856 ( .C1(n6604), .C2(n10365), .A(n6649), .B(n10364), .ZN(
        n10432) );
  OAI22_X1 U12857 ( .A1(n10367), .A2(n15069), .B1(n13868), .B2(n10366), .ZN(
        n10368) );
  AOI21_X1 U12858 ( .B1(n10432), .B2(n15064), .A(n10368), .ZN(n10373) );
  NAND2_X1 U12859 ( .A1(n10369), .A2(n12464), .ZN(n10371) );
  NAND2_X1 U12860 ( .A1(n6651), .A2(n13551), .ZN(n10370) );
  XNOR2_X1 U12861 ( .A(n10567), .B(n12466), .ZN(n10433) );
  NAND2_X1 U12862 ( .A1(n10433), .A2(n15072), .ZN(n10372) );
  OAI211_X1 U12863 ( .C1(n10374), .C2(n15075), .A(n10373), .B(n10372), .ZN(
        P2_U3253) );
  NAND2_X1 U12864 ( .A1(n10376), .A2(n10375), .ZN(n10377) );
  OR2_X1 U12865 ( .A1(n10379), .A2(n9924), .ZN(n10382) );
  AOI22_X1 U12866 ( .A1(n12116), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11366), 
        .B2(n10380), .ZN(n10381) );
  XNOR2_X1 U12867 ( .A(n14962), .B(n14258), .ZN(n12139) );
  XNOR2_X1 U12868 ( .A(n10546), .B(n10545), .ZN(n10397) );
  INV_X1 U12869 ( .A(n10397), .ZN(n14965) );
  NAND2_X1 U12870 ( .A1(n11381), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10390) );
  INV_X1 U12871 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10383) );
  AND2_X1 U12872 ( .A1(n10384), .A2(n10383), .ZN(n10385) );
  OR2_X1 U12873 ( .A1(n10385), .A2(n10536), .ZN(n14818) );
  OR2_X1 U12874 ( .A1(n6575), .A2(n14818), .ZN(n10389) );
  OR2_X1 U12875 ( .A1(n11919), .A2(n10386), .ZN(n10388) );
  OR2_X1 U12876 ( .A1(n9229), .A2(n8748), .ZN(n10387) );
  NAND4_X1 U12877 ( .A1(n10390), .A2(n10389), .A3(n10388), .A4(n10387), .ZN(
        n14257) );
  INV_X1 U12878 ( .A(n14257), .ZN(n14872) );
  OAI22_X1 U12879 ( .A1(n14869), .A2(n14517), .B1(n14872), .B2(n14637), .ZN(
        n10396) );
  OR2_X1 U12880 ( .A1(n14956), .A2(n14869), .ZN(n10391) );
  NAND2_X1 U12881 ( .A1(n10393), .A2(n10545), .ZN(n10394) );
  AOI21_X1 U12882 ( .B1(n10526), .B2(n10394), .A(n14724), .ZN(n10395) );
  AOI211_X1 U12883 ( .C1(n10397), .C2(n14729), .A(n10396), .B(n10395), .ZN(
        n14964) );
  MUX2_X1 U12884 ( .A(n10398), .B(n14964), .S(n14544), .Z(n10403) );
  AOI211_X1 U12885 ( .C1(n14962), .C2(n10399), .A(n14924), .B(n6800), .ZN(
        n14960) );
  INV_X1 U12886 ( .A(n14962), .ZN(n10400) );
  OAI22_X1 U12887 ( .A1(n10400), .A2(n14506), .B1(n14882), .B2(n14541), .ZN(
        n10401) );
  AOI21_X1 U12888 ( .B1(n14960), .B2(n14739), .A(n10401), .ZN(n10402) );
  OAI211_X1 U12889 ( .C1(n14965), .C2(n14508), .A(n10403), .B(n10402), .ZN(
        P1_U3284) );
  NAND2_X1 U12890 ( .A1(n10836), .A2(n12393), .ZN(n10405) );
  AOI22_X1 U12891 ( .A1(n11505), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n11504), 
        .B2(n15051), .ZN(n10404) );
  INV_X1 U12892 ( .A(n14017), .ZN(n10565) );
  INV_X1 U12893 ( .A(n10406), .ZN(n10408) );
  NAND2_X1 U12894 ( .A1(n10408), .A2(n10407), .ZN(n10409) );
  XNOR2_X1 U12895 ( .A(n14017), .B(n6627), .ZN(n11702) );
  AND2_X1 U12896 ( .A1(n13549), .A2(n6649), .ZN(n10411) );
  NAND2_X1 U12897 ( .A1(n11702), .A2(n10411), .ZN(n10713) );
  INV_X1 U12898 ( .A(n11702), .ZN(n10413) );
  INV_X1 U12899 ( .A(n10411), .ZN(n10412) );
  NAND2_X1 U12900 ( .A1(n10413), .A2(n10412), .ZN(n10414) );
  NAND2_X1 U12901 ( .A1(n10713), .A2(n10414), .ZN(n10415) );
  AOI21_X1 U12902 ( .B1(n10416), .B2(n10415), .A(n13478), .ZN(n10417) );
  NAND2_X1 U12903 ( .A1(n10417), .A2(n11704), .ZN(n10430) );
  NAND2_X1 U12904 ( .A1(n10418), .A2(n11706), .ZN(n10419) );
  NAND2_X1 U12905 ( .A1(n10654), .A2(n10419), .ZN(n10663) );
  NAND2_X1 U12906 ( .A1(n11619), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n10421) );
  NAND2_X1 U12907 ( .A1(n11618), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n10420) );
  AND2_X1 U12908 ( .A1(n10421), .A2(n10420), .ZN(n10423) );
  NAND2_X1 U12909 ( .A1(n12390), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n10422) );
  OAI211_X1 U12910 ( .C1(n10663), .C2(n11606), .A(n10423), .B(n10422), .ZN(
        n13548) );
  NAND2_X1 U12911 ( .A1(n13548), .A2(n13517), .ZN(n10425) );
  NAND2_X1 U12912 ( .A1(n13550), .A2(n13518), .ZN(n10424) );
  NAND2_X1 U12913 ( .A1(n10425), .A2(n10424), .ZN(n10560) );
  INV_X1 U12914 ( .A(n10560), .ZN(n10427) );
  OAI22_X1 U12915 ( .A1(n13503), .A2(n10427), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10426), .ZN(n10428) );
  AOI21_X1 U12916 ( .B1(n10563), .B2(n13522), .A(n10428), .ZN(n10429) );
  OAI211_X1 U12917 ( .C1(n10565), .C2(n13525), .A(n10430), .B(n10429), .ZN(
        P2_U3206) );
  AOI211_X1 U12918 ( .C1(n14012), .C2(n10433), .A(n10432), .B(n10431), .ZN(
        n10436) );
  AOI22_X1 U12919 ( .A1(n6604), .A2(n14051), .B1(P2_REG0_REG_12__SCAN_IN), 
        .B2(n15104), .ZN(n10434) );
  OAI21_X1 U12920 ( .B1(n10436), .B2(n15104), .A(n10434), .ZN(P2_U3466) );
  AOI22_X1 U12921 ( .A1(n6604), .A2(n13992), .B1(P2_REG1_REG_12__SCAN_IN), 
        .B2(n15109), .ZN(n10435) );
  OAI21_X1 U12922 ( .B1(n10436), .B2(n15109), .A(n10435), .ZN(P2_U3511) );
  OAI22_X1 U12923 ( .A1(n15165), .A2(n12787), .B1(n10437), .B2(n15169), .ZN(
        n10440) );
  MUX2_X1 U12924 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n10438), .S(n15204), .Z(
        n10439) );
  AOI211_X1 U12925 ( .C1(n13270), .C2(n10441), .A(n10440), .B(n10439), .ZN(
        n10442) );
  INV_X1 U12926 ( .A(n10442), .ZN(P3_U3229) );
  MUX2_X1 U12927 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n11907), .Z(n10740) );
  XNOR2_X1 U12928 ( .A(n10742), .B(n10741), .ZN(n11525) );
  INV_X1 U12929 ( .A(n11525), .ZN(n10445) );
  OAI222_X1 U12930 ( .A1(P2_U3088), .A2(n12179), .B1(n14088), .B2(n10445), 
        .C1(n13615), .C2(n14086), .ZN(P2_U3306) );
  OAI222_X1 U12931 ( .A1(n11931), .A2(P1_U3086), .B1(n14694), .B2(n10445), 
        .C1(n13655), .C2(n14684), .ZN(P1_U3334) );
  OAI21_X1 U12932 ( .B1(n10447), .B2(n12928), .A(n10446), .ZN(n10646) );
  NAND2_X1 U12933 ( .A1(n10578), .A2(n10448), .ZN(n10599) );
  NAND2_X1 U12934 ( .A1(n10578), .A2(n10449), .ZN(n10450) );
  NAND2_X1 U12935 ( .A1(n10450), .A2(n12928), .ZN(n10451) );
  NAND3_X1 U12936 ( .A1(n10599), .A2(n14762), .A3(n10451), .ZN(n10453) );
  AOI22_X1 U12937 ( .A1(n15195), .A2(n12972), .B1(n12974), .B2(n15192), .ZN(
        n10452) );
  NAND2_X1 U12938 ( .A1(n10453), .A2(n10452), .ZN(n10643) );
  AOI21_X1 U12939 ( .B1(n14798), .B2(n10646), .A(n10643), .ZN(n10501) );
  INV_X1 U12940 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n10454) );
  OAI22_X1 U12941 ( .A1(n10642), .A2(n13384), .B1(n15232), .B2(n10454), .ZN(
        n10455) );
  INV_X1 U12942 ( .A(n10455), .ZN(n10456) );
  OAI21_X1 U12943 ( .B1(n10501), .B2(n15234), .A(n10456), .ZN(P3_U3408) );
  INV_X1 U12944 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10914) );
  NOR2_X1 U12945 ( .A1(n10914), .A2(n10458), .ZN(n10625) );
  AOI211_X1 U12946 ( .C1(n10458), .C2(n10914), .A(n10625), .B(n15046), .ZN(
        n10459) );
  INV_X1 U12947 ( .A(n10459), .ZN(n10471) );
  INV_X1 U12948 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10721) );
  NOR2_X1 U12949 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10721), .ZN(n10469) );
  OR2_X1 U12950 ( .A1(n10461), .A2(n10460), .ZN(n10464) );
  INV_X1 U12951 ( .A(n10462), .ZN(n10463) );
  INV_X1 U12952 ( .A(n10629), .ZN(n10465) );
  XNOR2_X1 U12953 ( .A(n10682), .B(n10465), .ZN(n10466) );
  NAND2_X1 U12954 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n10466), .ZN(n10630) );
  OAI211_X1 U12955 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n10466), .A(n15039), 
        .B(n10630), .ZN(n10467) );
  INV_X1 U12956 ( .A(n10467), .ZN(n10468) );
  AOI211_X1 U12957 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n14987), .A(n10469), 
        .B(n10468), .ZN(n10470) );
  OAI211_X1 U12958 ( .C1(n14993), .C2(n10623), .A(n10471), .B(n10470), .ZN(
        P2_U3229) );
  OR2_X1 U12959 ( .A1(n10969), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n10473) );
  NAND2_X1 U12960 ( .A1(n10473), .A2(n10472), .ZN(n10474) );
  INV_X1 U12961 ( .A(n10474), .ZN(n10475) );
  XNOR2_X1 U12962 ( .A(n10474), .B(n14902), .ZN(n14899) );
  INV_X1 U12963 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14898) );
  NAND2_X1 U12964 ( .A1(n14899), .A2(n14898), .ZN(n14897) );
  OAI21_X1 U12965 ( .B1(n10475), .B2(n14902), .A(n14897), .ZN(n10477) );
  INV_X1 U12966 ( .A(n11054), .ZN(n11169) );
  XNOR2_X1 U12967 ( .A(n11169), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n10476) );
  NOR2_X1 U12968 ( .A1(n10477), .A2(n10476), .ZN(n11048) );
  AOI211_X1 U12969 ( .C1(n10477), .C2(n10476), .A(n11048), .B(n14323), .ZN(
        n10490) );
  NAND2_X1 U12970 ( .A1(n10969), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10479) );
  NAND2_X1 U12971 ( .A1(n10479), .A2(n10478), .ZN(n10480) );
  INV_X1 U12972 ( .A(n10480), .ZN(n10482) );
  XNOR2_X1 U12973 ( .A(n10480), .B(n14902), .ZN(n14896) );
  NOR2_X1 U12974 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14896), .ZN(n14895) );
  AOI21_X1 U12975 ( .B1(n10482), .B2(n10481), .A(n14895), .ZN(n10485) );
  INV_X1 U12976 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10483) );
  MUX2_X1 U12977 ( .A(n10483), .B(P1_REG2_REG_16__SCAN_IN), .S(n11054), .Z(
        n10484) );
  NAND2_X1 U12978 ( .A1(n10484), .A2(n10485), .ZN(n11053) );
  OAI211_X1 U12979 ( .C1(n10485), .C2(n10484), .A(n14318), .B(n11053), .ZN(
        n10488) );
  INV_X1 U12980 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n13714) );
  NOR2_X1 U12981 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13714), .ZN(n10486) );
  AOI21_X1 U12982 ( .B1(n14891), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10486), 
        .ZN(n10487) );
  OAI211_X1 U12983 ( .C1(n14320), .C2(n11054), .A(n10488), .B(n10487), .ZN(
        n10489) );
  OR2_X1 U12984 ( .A1(n10490), .A2(n10489), .ZN(P1_U3259) );
  INV_X1 U12985 ( .A(n13334), .ZN(n10499) );
  AOI22_X1 U12986 ( .A1(n10499), .A2(n10491), .B1(n15241), .B2(
        P3_REG1_REG_4__SCAN_IN), .ZN(n10492) );
  OAI21_X1 U12987 ( .B1(n10493), .B2(n15241), .A(n10492), .ZN(P3_U3463) );
  INV_X1 U12988 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10494) );
  OAI22_X1 U12989 ( .A1(n13334), .A2(n10495), .B1(n15240), .B2(n10494), .ZN(
        n10496) );
  AOI21_X1 U12990 ( .B1(n10497), .B2(n15240), .A(n10496), .ZN(n10498) );
  INV_X1 U12991 ( .A(n10498), .ZN(P3_U3462) );
  AOI22_X1 U12992 ( .A1(n10499), .A2(n10669), .B1(n15241), .B2(
        P3_REG1_REG_6__SCAN_IN), .ZN(n10500) );
  OAI21_X1 U12993 ( .B1(n10501), .B2(n15241), .A(n10500), .ZN(P3_U3465) );
  MUX2_X1 U12994 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13037), .Z(n10765) );
  XNOR2_X1 U12995 ( .A(n10765), .B(n10767), .ZN(n10768) );
  XOR2_X1 U12996 ( .A(n10768), .B(n10769), .Z(n10518) );
  NAND2_X1 U12997 ( .A1(n10508), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n10506) );
  NAND2_X1 U12998 ( .A1(n10506), .A2(n10505), .ZN(n10788) );
  XNOR2_X1 U12999 ( .A(n10788), .B(n10767), .ZN(n10507) );
  NAND2_X1 U13000 ( .A1(P3_REG2_REG_11__SCAN_IN), .A2(n10507), .ZN(n10790) );
  OAI21_X1 U13001 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n10507), .A(n10790), 
        .ZN(n10516) );
  AND2_X1 U13002 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n12703) );
  AOI21_X1 U13003 ( .B1(n15113), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n12703), 
        .ZN(n10514) );
  NAND2_X1 U13004 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n10508), .ZN(n10510) );
  NAND2_X1 U13005 ( .A1(n10510), .A2(n10509), .ZN(n10774) );
  XNOR2_X1 U13006 ( .A(n10767), .B(n10774), .ZN(n10511) );
  NAND2_X1 U13007 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n10511), .ZN(n10775) );
  OAI21_X1 U13008 ( .B1(n10511), .B2(P3_REG1_REG_11__SCAN_IN), .A(n10775), 
        .ZN(n10512) );
  NAND2_X1 U13009 ( .A1(n13023), .A2(n10512), .ZN(n10513) );
  OAI211_X1 U13010 ( .C1(n15150), .C2(n10789), .A(n10514), .B(n10513), .ZN(
        n10515) );
  AOI21_X1 U13011 ( .B1(n10516), .B2(n15154), .A(n10515), .ZN(n10517) );
  OAI21_X1 U13012 ( .B1(n10518), .B2(n13078), .A(n10517), .ZN(P3_U3193) );
  NAND2_X1 U13013 ( .A1(n11459), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10524) );
  INV_X1 U13014 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10519) );
  OR2_X1 U13015 ( .A1(n11921), .A2(n10519), .ZN(n10523) );
  OR2_X1 U13016 ( .A1(n10538), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10520) );
  NAND2_X1 U13017 ( .A1(n10841), .A2(n10520), .ZN(n14730) );
  OR2_X1 U13018 ( .A1(n6575), .A2(n14730), .ZN(n10522) );
  OR2_X1 U13019 ( .A1(n11919), .A2(n14750), .ZN(n10521) );
  NAND4_X1 U13020 ( .A1(n10524), .A2(n10523), .A3(n10522), .A4(n10521), .ZN(
        n14255) );
  INV_X1 U13021 ( .A(n14255), .ZN(n14819) );
  NAND2_X1 U13022 ( .A1(n14962), .A2(n14807), .ZN(n10525) );
  AOI22_X1 U13023 ( .A1(n12116), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n11366), 
        .B2(n10528), .ZN(n10529) );
  XNOR2_X1 U13024 ( .A(n14806), .B(n14257), .ZN(n12140) );
  OR2_X1 U13025 ( .A1(n14806), .A2(n14872), .ZN(n10531) );
  NAND2_X1 U13026 ( .A1(n10532), .A2(n11913), .ZN(n10535) );
  AOI22_X1 U13027 ( .A1(n12116), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n11366), 
        .B2(n10533), .ZN(n10534) );
  NAND2_X1 U13028 ( .A1(n11381), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10543) );
  NOR2_X1 U13029 ( .A1(n10536), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10537) );
  OR2_X1 U13030 ( .A1(n10538), .A2(n10537), .ZN(n14831) );
  OR2_X1 U13031 ( .A1(n6575), .A2(n14831), .ZN(n10542) );
  OR2_X1 U13032 ( .A1(n11919), .A2(n10539), .ZN(n10541) );
  OR2_X1 U13033 ( .A1(n9229), .A2(n9051), .ZN(n10540) );
  NAND4_X1 U13034 ( .A1(n10543), .A2(n10542), .A3(n10541), .A4(n10540), .ZN(
        n14256) );
  XNOR2_X1 U13035 ( .A(n14828), .B(n14256), .ZN(n12142) );
  XNOR2_X1 U13036 ( .A(n10851), .B(n12142), .ZN(n10544) );
  OAI222_X1 U13037 ( .A1(n14637), .A2(n14819), .B1(n10544), .B2(n14724), .C1(
        n14517), .C2(n14872), .ZN(n10758) );
  INV_X1 U13038 ( .A(n10758), .ZN(n10556) );
  OR2_X1 U13039 ( .A1(n14962), .A2(n14258), .ZN(n10547) );
  NOR2_X1 U13040 ( .A1(n14806), .A2(n14257), .ZN(n10548) );
  XNOR2_X1 U13041 ( .A(n10829), .B(n12142), .ZN(n10760) );
  INV_X1 U13042 ( .A(n14546), .ZN(n14474) );
  AND2_X1 U13043 ( .A1(n14828), .A2(n10705), .ZN(n10549) );
  OR2_X1 U13044 ( .A1(n10549), .A2(n14737), .ZN(n10757) );
  NAND2_X1 U13045 ( .A1(n14743), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10550) );
  OAI21_X1 U13046 ( .B1(n14541), .B2(n14831), .A(n10550), .ZN(n10551) );
  AOI21_X1 U13047 ( .B1(n14828), .B2(n14733), .A(n10551), .ZN(n10552) );
  OAI21_X1 U13048 ( .B1(n10757), .B2(n10553), .A(n10552), .ZN(n10554) );
  AOI21_X1 U13049 ( .B1(n10760), .B2(n14474), .A(n10554), .ZN(n10555) );
  OAI21_X1 U13050 ( .B1(n10556), .B2(n14743), .A(n10555), .ZN(P1_U3282) );
  INV_X1 U13051 ( .A(n13550), .ZN(n10557) );
  OR2_X1 U13052 ( .A1(n6604), .A2(n10557), .ZN(n10558) );
  XNOR2_X1 U13053 ( .A(n14017), .B(n13549), .ZN(n12465) );
  INV_X1 U13054 ( .A(n12465), .ZN(n10569) );
  OAI21_X1 U13055 ( .B1(n6543), .B2(n12465), .A(n10652), .ZN(n10561) );
  AOI21_X1 U13056 ( .B1(n10561), .B2(n13891), .A(n10560), .ZN(n14019) );
  AOI211_X1 U13057 ( .C1(n14017), .C2(n10562), .A(n6649), .B(n6955), .ZN(
        n14016) );
  AOI22_X1 U13058 ( .A1(n15075), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n10563), 
        .B2(n15062), .ZN(n10564) );
  OAI21_X1 U13059 ( .B1(n10565), .B2(n15069), .A(n10564), .ZN(n10571) );
  NAND2_X1 U13060 ( .A1(n6604), .A2(n13550), .ZN(n10568) );
  XNOR2_X1 U13061 ( .A(n10661), .B(n10569), .ZN(n14020) );
  NOR2_X1 U13062 ( .A1(n14020), .A2(n13871), .ZN(n10570) );
  AOI211_X1 U13063 ( .C1(n14016), .C2(n15064), .A(n10571), .B(n10570), .ZN(
        n10572) );
  OAI21_X1 U13064 ( .B1(n15075), .B2(n14019), .A(n10572), .ZN(P2_U3252) );
  INV_X1 U13065 ( .A(n12931), .ZN(n10573) );
  XNOR2_X1 U13066 ( .A(n10574), .B(n10573), .ZN(n15215) );
  INV_X1 U13067 ( .A(n15183), .ZN(n10575) );
  NAND2_X1 U13068 ( .A1(n15204), .A2(n10575), .ZN(n13116) );
  NAND2_X1 U13069 ( .A1(n10576), .A2(n12931), .ZN(n10577) );
  NAND2_X1 U13070 ( .A1(n10578), .A2(n10577), .ZN(n10579) );
  NAND2_X1 U13071 ( .A1(n10579), .A2(n14762), .ZN(n10581) );
  AOI22_X1 U13072 ( .A1(n15192), .A2(n12975), .B1(n12973), .B2(n15195), .ZN(
        n10580) );
  OAI211_X1 U13073 ( .C1(n15177), .C2(n15215), .A(n10581), .B(n10580), .ZN(
        n15216) );
  MUX2_X1 U13074 ( .A(n15216), .B(P3_REG2_REG_5__SCAN_IN), .S(n15206), .Z(
        n10582) );
  INV_X1 U13075 ( .A(n10582), .ZN(n10586) );
  NOR2_X1 U13076 ( .A1(n10583), .A2(n15226), .ZN(n15217) );
  AOI22_X1 U13077 ( .A1(n14770), .A2(n15217), .B1(n15201), .B2(n10584), .ZN(
        n10585) );
  OAI211_X1 U13078 ( .C1(n15215), .C2(n13116), .A(n10586), .B(n10585), .ZN(
        P3_U3228) );
  INV_X1 U13079 ( .A(n10587), .ZN(n10595) );
  NAND2_X1 U13080 ( .A1(n10588), .A2(n15064), .ZN(n10591) );
  AOI22_X1 U13081 ( .A1(n15075), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n10589), 
        .B2(n15062), .ZN(n10590) );
  OAI211_X1 U13082 ( .C1(n6950), .C2(n15069), .A(n10591), .B(n10590), .ZN(
        n10592) );
  AOI21_X1 U13083 ( .B1(n10593), .B2(n13868), .A(n10592), .ZN(n10594) );
  OAI21_X1 U13084 ( .B1(n10595), .B2(n13871), .A(n10594), .ZN(P2_U3255) );
  OAI21_X1 U13085 ( .B1(n10597), .B2(n7795), .A(n10596), .ZN(n10755) );
  NAND2_X1 U13086 ( .A1(n10599), .A2(n10598), .ZN(n10600) );
  OAI211_X1 U13087 ( .C1(n10600), .C2(n12933), .A(n10814), .B(n14762), .ZN(
        n10602) );
  AOI22_X1 U13088 ( .A1(n15192), .A2(n12973), .B1(n12971), .B2(n15195), .ZN(
        n10601) );
  NAND2_X1 U13089 ( .A1(n10602), .A2(n10601), .ZN(n10752) );
  AOI21_X1 U13090 ( .B1(n14798), .B2(n10755), .A(n10752), .ZN(n10608) );
  OAI22_X1 U13091 ( .A1(n13334), .A2(n12806), .B1(n15240), .B2(n9982), .ZN(
        n10603) );
  INV_X1 U13092 ( .A(n10603), .ZN(n10604) );
  OAI21_X1 U13093 ( .B1(n10608), .B2(n15241), .A(n10604), .ZN(P3_U3466) );
  INV_X1 U13094 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n10605) );
  OAI22_X1 U13095 ( .A1(n12806), .A2(n13384), .B1(n15232), .B2(n10605), .ZN(
        n10606) );
  INV_X1 U13096 ( .A(n10606), .ZN(n10607) );
  OAI21_X1 U13097 ( .B1(n10608), .B2(n15234), .A(n10607), .ZN(P3_U3411) );
  INV_X1 U13098 ( .A(n10609), .ZN(n10751) );
  OR2_X1 U13099 ( .A1(n10612), .A2(n12974), .ZN(n10613) );
  XNOR2_X1 U13100 ( .A(n12614), .B(n10669), .ZN(n10614) );
  XOR2_X1 U13101 ( .A(n12973), .B(n10614), .Z(n10674) );
  INV_X1 U13102 ( .A(n10614), .ZN(n10615) );
  NAND2_X1 U13103 ( .A1(n10615), .A2(n12973), .ZN(n10616) );
  NAND2_X1 U13104 ( .A1(n10671), .A2(n10616), .ZN(n10617) );
  XNOR2_X1 U13105 ( .A(n12933), .B(n12548), .ZN(n10728) );
  OAI211_X1 U13106 ( .C1(n10617), .C2(n10728), .A(n10731), .B(n12673), .ZN(
        n10622) );
  OAI22_X1 U13107 ( .A1(n12720), .A2(n12806), .B1(n10618), .B2(n12719), .ZN(
        n10619) );
  AOI211_X1 U13108 ( .C1(n12717), .C2(n12971), .A(n10620), .B(n10619), .ZN(
        n10621) );
  OAI211_X1 U13109 ( .C1(n10751), .C2(n12706), .A(n10622), .B(n10621), .ZN(
        P3_U3153) );
  NOR2_X1 U13110 ( .A1(n10624), .A2(n10623), .ZN(n10626) );
  XNOR2_X1 U13111 ( .A(n10923), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n10627) );
  NOR2_X1 U13112 ( .A1(n10628), .A2(n10627), .ZN(n10894) );
  AOI211_X1 U13113 ( .C1(n10628), .C2(n10627), .A(n15046), .B(n10894), .ZN(
        n10640) );
  NAND2_X1 U13114 ( .A1(n10682), .A2(n10629), .ZN(n10631) );
  NAND2_X1 U13115 ( .A1(n10923), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n10898) );
  OAI21_X1 U13116 ( .B1(n10923), .B2(P2_REG2_REG_16__SCAN_IN), .A(n10898), 
        .ZN(n10632) );
  INV_X1 U13117 ( .A(n10632), .ZN(n10633) );
  NAND2_X1 U13118 ( .A1(n10634), .A2(n10633), .ZN(n10899) );
  OAI211_X1 U13119 ( .C1(n10634), .C2(n10633), .A(n10899), .B(n15039), .ZN(
        n10637) );
  INV_X1 U13120 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n11109) );
  NOR2_X1 U13121 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11109), .ZN(n10635) );
  AOI21_X1 U13122 ( .B1(n14987), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n10635), 
        .ZN(n10636) );
  OAI211_X1 U13123 ( .C1(n14993), .C2(n10638), .A(n10637), .B(n10636), .ZN(
        n10639) );
  OR2_X1 U13124 ( .A1(n10640), .A2(n10639), .ZN(P2_U3230) );
  INV_X1 U13125 ( .A(n10677), .ZN(n10641) );
  OAI22_X1 U13126 ( .A1(n15165), .A2(n10642), .B1(n10641), .B2(n15169), .ZN(
        n10645) );
  MUX2_X1 U13127 ( .A(n10643), .B(P3_REG2_REG_6__SCAN_IN), .S(n15206), .Z(
        n10644) );
  AOI211_X1 U13128 ( .C1(n13270), .C2(n10646), .A(n10645), .B(n10644), .ZN(
        n10647) );
  INV_X1 U13129 ( .A(n10647), .ZN(P3_U3227) );
  NAND2_X1 U13130 ( .A1(n10968), .A2(n12393), .ZN(n10650) );
  AOI22_X1 U13131 ( .A1(n11505), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n11504), 
        .B2(n10648), .ZN(n10649) );
  XNOR2_X1 U13132 ( .A(n6593), .B(n13548), .ZN(n12468) );
  INV_X1 U13133 ( .A(n13549), .ZN(n12290) );
  NAND2_X1 U13134 ( .A1(n14017), .A2(n12290), .ZN(n10651) );
  XOR2_X1 U13135 ( .A(n12468), .B(n10681), .Z(n10659) );
  INV_X1 U13136 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n10917) );
  NAND2_X1 U13137 ( .A1(n10654), .A2(n10721), .ZN(n10655) );
  NAND2_X1 U13138 ( .A1(n10686), .A2(n10655), .ZN(n10720) );
  OR2_X1 U13139 ( .A1(n10720), .A2(n11606), .ZN(n10657) );
  AOI22_X1 U13140 ( .A1(n12390), .A2(P2_REG1_REG_15__SCAN_IN), .B1(n10688), 
        .B2(P2_REG2_REG_15__SCAN_IN), .ZN(n10656) );
  OAI211_X1 U13141 ( .C1(n8942), .C2(n10917), .A(n10657), .B(n10656), .ZN(
        n13547) );
  AND2_X1 U13142 ( .A1(n13549), .A2(n13518), .ZN(n10658) );
  AOI21_X1 U13143 ( .B1(n13547), .B2(n13517), .A(n10658), .ZN(n11707) );
  OAI21_X1 U13144 ( .B1(n10659), .B2(n13875), .A(n11707), .ZN(n10872) );
  INV_X1 U13145 ( .A(n10872), .ZN(n10668) );
  AND2_X1 U13146 ( .A1(n14017), .A2(n13549), .ZN(n10660) );
  XOR2_X1 U13147 ( .A(n12468), .B(n10698), .Z(n10874) );
  AOI211_X1 U13148 ( .C1(n6593), .C2(n10662), .A(n6649), .B(n10694), .ZN(
        n10873) );
  NAND2_X1 U13149 ( .A1(n10873), .A2(n15064), .ZN(n10665) );
  INV_X1 U13150 ( .A(n10663), .ZN(n11709) );
  AOI22_X1 U13151 ( .A1(n15075), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11709), 
        .B2(n15062), .ZN(n10664) );
  OAI211_X1 U13152 ( .C1(n6959), .C2(n15069), .A(n10665), .B(n10664), .ZN(
        n10666) );
  AOI21_X1 U13153 ( .B1(n10874), .B2(n15072), .A(n10666), .ZN(n10667) );
  OAI21_X1 U13154 ( .B1(n10668), .B2(n15075), .A(n10667), .ZN(P2_U3251) );
  AOI22_X1 U13155 ( .A1(n12737), .A2(n10669), .B1(n12731), .B2(n12974), .ZN(
        n10670) );
  NAND2_X1 U13156 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n15131) );
  OAI211_X1 U13157 ( .C1(n12805), .C2(n12734), .A(n10670), .B(n15131), .ZN(
        n10676) );
  INV_X1 U13158 ( .A(n10671), .ZN(n10672) );
  AOI211_X1 U13159 ( .C1(n10674), .C2(n10673), .A(n12739), .B(n10672), .ZN(
        n10675) );
  AOI211_X1 U13160 ( .C1(n10677), .C2(n12729), .A(n10676), .B(n10675), .ZN(
        n10678) );
  INV_X1 U13161 ( .A(n10678), .ZN(P3_U3179) );
  INV_X1 U13162 ( .A(n10720), .ZN(n10693) );
  INV_X1 U13163 ( .A(n13548), .ZN(n10679) );
  AND2_X1 U13164 ( .A1(n6593), .A2(n10679), .ZN(n10680) );
  NAND2_X1 U13165 ( .A1(n11178), .A2(n12393), .ZN(n10684) );
  AOI22_X1 U13166 ( .A1(n11505), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n11504), 
        .B2(n10682), .ZN(n10683) );
  INV_X1 U13167 ( .A(n13547), .ZN(n10929) );
  XNOR2_X1 U13168 ( .A(n12300), .B(n10929), .ZN(n12470) );
  INV_X1 U13169 ( .A(n12470), .ZN(n10920) );
  XNOR2_X1 U13170 ( .A(n10928), .B(n10920), .ZN(n10692) );
  INV_X1 U13171 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n10691) );
  INV_X1 U13172 ( .A(n10686), .ZN(n10685) );
  NAND2_X1 U13173 ( .A1(n10686), .A2(n11109), .ZN(n10687) );
  NAND2_X1 U13174 ( .A1(n10934), .A2(n10687), .ZN(n11108) );
  OR2_X1 U13175 ( .A1(n11108), .A2(n11606), .ZN(n10690) );
  AOI22_X1 U13176 ( .A1(n11619), .A2(P2_REG0_REG_16__SCAN_IN), .B1(n10688), 
        .B2(P2_REG2_REG_16__SCAN_IN), .ZN(n10689) );
  OAI211_X1 U13177 ( .C1(n11609), .C2(n10691), .A(n10690), .B(n10689), .ZN(
        n13546) );
  AOI22_X1 U13178 ( .A1(n13546), .A2(n13517), .B1(n13518), .B2(n13548), .ZN(
        n10722) );
  OAI21_X1 U13179 ( .B1(n10692), .B2(n13875), .A(n10722), .ZN(n10911) );
  AOI21_X1 U13180 ( .B1(n10693), .B2(n15062), .A(n10911), .ZN(n10703) );
  INV_X1 U13181 ( .A(n10694), .ZN(n10695) );
  AOI211_X1 U13182 ( .C1(n12300), .C2(n10695), .A(n6649), .B(n10943), .ZN(
        n10912) );
  INV_X1 U13183 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n10696) );
  OAI22_X1 U13184 ( .A1(n10919), .A2(n15069), .B1(n13868), .B2(n10696), .ZN(
        n10697) );
  AOI21_X1 U13185 ( .B1(n10912), .B2(n15064), .A(n10697), .ZN(n10702) );
  NAND2_X1 U13186 ( .A1(n6593), .A2(n13548), .ZN(n10699) );
  XNOR2_X1 U13187 ( .A(n10921), .B(n10920), .ZN(n10913) );
  NAND2_X1 U13188 ( .A1(n10913), .A2(n15072), .ZN(n10701) );
  OAI211_X1 U13189 ( .C1(n10703), .C2(n15075), .A(n10702), .B(n10701), .ZN(
        P2_U3250) );
  XNOR2_X1 U13190 ( .A(n10704), .B(n12140), .ZN(n14970) );
  INV_X1 U13191 ( .A(n14256), .ZN(n14808) );
  OAI211_X1 U13192 ( .C1(n6799), .C2(n6800), .A(n14736), .B(n10705), .ZN(
        n10706) );
  OAI21_X1 U13193 ( .B1(n14808), .B2(n14637), .A(n10706), .ZN(n14971) );
  OAI22_X1 U13194 ( .A1(n6799), .A2(n14506), .B1(n14541), .B2(n14818), .ZN(
        n10711) );
  OAI211_X1 U13195 ( .C1(n10708), .C2(n12140), .A(n10707), .B(n14832), .ZN(
        n10709) );
  OAI21_X1 U13196 ( .B1(n14807), .B2(n14517), .A(n10709), .ZN(n14973) );
  MUX2_X1 U13197 ( .A(n14973), .B(P1_REG2_REG_10__SCAN_IN), .S(n14743), .Z(
        n10710) );
  AOI211_X1 U13198 ( .C1(n14739), .C2(n14971), .A(n10711), .B(n10710), .ZN(
        n10712) );
  OAI21_X1 U13199 ( .B1(n14546), .B2(n14970), .A(n10712), .ZN(P1_U3283) );
  XNOR2_X1 U13200 ( .A(n12294), .B(n6627), .ZN(n10714) );
  NAND2_X1 U13201 ( .A1(n13548), .A2(n13845), .ZN(n10715) );
  XNOR2_X1 U13202 ( .A(n10714), .B(n10715), .ZN(n11705) );
  INV_X1 U13203 ( .A(n10714), .ZN(n10716) );
  NAND2_X1 U13204 ( .A1(n10716), .A2(n10715), .ZN(n10717) );
  XNOR2_X1 U13205 ( .A(n12300), .B(n6627), .ZN(n11064) );
  AOI22_X1 U13206 ( .A1(n10719), .A2(n13527), .B1(n13436), .B2(n13547), .ZN(
        n10727) );
  AND2_X1 U13207 ( .A1(n13547), .A2(n6649), .ZN(n10718) );
  INV_X1 U13208 ( .A(n6564), .ZN(n10726) );
  NOR2_X1 U13209 ( .A1(n13495), .A2(n10720), .ZN(n10724) );
  OAI22_X1 U13210 ( .A1(n13503), .A2(n10722), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10721), .ZN(n10723) );
  AOI211_X1 U13211 ( .C1(n12300), .C2(n13510), .A(n10724), .B(n10723), .ZN(
        n10725) );
  OAI21_X1 U13212 ( .B1(n10727), .B2(n10726), .A(n10725), .ZN(P2_U3213) );
  INV_X1 U13213 ( .A(n10823), .ZN(n10739) );
  INV_X1 U13214 ( .A(n10728), .ZN(n10729) );
  NAND2_X1 U13215 ( .A1(n10729), .A2(n12972), .ZN(n10730) );
  XNOR2_X1 U13216 ( .A(n12614), .B(n10732), .ZN(n10951) );
  XNOR2_X1 U13217 ( .A(n10951), .B(n12971), .ZN(n10733) );
  NAND2_X1 U13218 ( .A1(n10734), .A2(n10733), .ZN(n10954) );
  OAI211_X1 U13219 ( .C1(n10734), .C2(n10733), .A(n10954), .B(n12673), .ZN(
        n10738) );
  NAND2_X1 U13220 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n15155) );
  INV_X1 U13221 ( .A(n15155), .ZN(n10736) );
  OAI22_X1 U13222 ( .A1(n12720), .A2(n10822), .B1(n12805), .B2(n12719), .ZN(
        n10735) );
  AOI211_X1 U13223 ( .C1(n12717), .C2(n12970), .A(n10736), .B(n10735), .ZN(
        n10737) );
  OAI211_X1 U13224 ( .C1(n10739), .C2(n12706), .A(n10738), .B(n10737), .ZN(
        P3_U3161) );
  INV_X1 U13225 ( .A(SI_22_), .ZN(n10743) );
  NAND2_X1 U13226 ( .A1(n10744), .A2(n10743), .ZN(n10745) );
  MUX2_X1 U13227 ( .A(n10746), .B(n11538), .S(n11907), .Z(n10747) );
  NAND2_X1 U13228 ( .A1(n11402), .A2(n10747), .ZN(n10748) );
  AND2_X1 U13229 ( .A1(n10799), .A2(n10748), .ZN(n11537) );
  INV_X1 U13230 ( .A(n11537), .ZN(n10749) );
  OAI222_X1 U13231 ( .A1(n14086), .A2(n11538), .B1(P2_U3088), .B2(n6667), .C1(
        n14088), .C2(n10749), .ZN(P2_U3305) );
  OAI22_X1 U13232 ( .A1(n15165), .A2(n12806), .B1(n10751), .B2(n15169), .ZN(
        n10754) );
  MUX2_X1 U13233 ( .A(n10752), .B(P3_REG2_REG_7__SCAN_IN), .S(n15206), .Z(
        n10753) );
  AOI211_X1 U13234 ( .C1(n13270), .C2(n10755), .A(n10754), .B(n10753), .ZN(
        n10756) );
  INV_X1 U13235 ( .A(n10756), .ZN(P3_U3226) );
  INV_X1 U13236 ( .A(n14828), .ZN(n10849) );
  OAI22_X1 U13237 ( .A1(n10757), .A2(n14924), .B1(n10849), .B2(n14949), .ZN(
        n10759) );
  AOI211_X1 U13238 ( .C1(n14927), .C2(n10760), .A(n10759), .B(n10758), .ZN(
        n10762) );
  OR2_X1 U13239 ( .A1(n10762), .A2(n14984), .ZN(n10761) );
  OAI21_X1 U13240 ( .B1(n14986), .B2(n10539), .A(n10761), .ZN(P1_U3539) );
  INV_X1 U13241 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10764) );
  OR2_X1 U13242 ( .A1(n10762), .A2(n14975), .ZN(n10763) );
  OAI21_X1 U13243 ( .B1(n14953), .B2(n10764), .A(n10763), .ZN(P1_U3492) );
  MUX2_X1 U13244 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13037), .Z(n11118) );
  XNOR2_X1 U13245 ( .A(n11118), .B(n11127), .ZN(n10773) );
  INV_X1 U13246 ( .A(n12985), .ZN(n10778) );
  MUX2_X1 U13247 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13037), .Z(n10770) );
  INV_X1 U13248 ( .A(n10770), .ZN(n10771) );
  INV_X1 U13249 ( .A(n10765), .ZN(n10766) );
  XOR2_X1 U13250 ( .A(n12985), .B(n10770), .Z(n12978) );
  NAND2_X1 U13251 ( .A1(n12979), .A2(n12978), .ZN(n12977) );
  OAI21_X1 U13252 ( .B1(n10778), .B2(n10771), .A(n12977), .ZN(n10772) );
  NOR2_X1 U13253 ( .A1(n10772), .A2(n10773), .ZN(n11119) );
  AOI21_X1 U13254 ( .B1(n10773), .B2(n10772), .A(n11119), .ZN(n10797) );
  INV_X1 U13255 ( .A(n11127), .ZN(n11121) );
  INV_X1 U13256 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n10784) );
  NAND2_X1 U13257 ( .A1(n12985), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n10779) );
  NAND2_X1 U13258 ( .A1(n10789), .A2(n10774), .ZN(n10776) );
  NAND2_X1 U13259 ( .A1(n10776), .A2(n10775), .ZN(n12981) );
  INV_X1 U13260 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14794) );
  INV_X1 U13261 ( .A(n10779), .ZN(n10777) );
  AOI21_X1 U13262 ( .B1(n10778), .B2(n14794), .A(n10777), .ZN(n12982) );
  NAND2_X1 U13263 ( .A1(n12981), .A2(n12982), .ZN(n12980) );
  NAND2_X1 U13264 ( .A1(n10779), .A2(n12980), .ZN(n11126) );
  XNOR2_X1 U13265 ( .A(n11121), .B(n11126), .ZN(n10780) );
  NAND2_X1 U13266 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n10780), .ZN(n11128) );
  OAI21_X1 U13267 ( .B1(n10780), .B2(P3_REG1_REG_13__SCAN_IN), .A(n11128), 
        .ZN(n10781) );
  NAND2_X1 U13268 ( .A1(n13023), .A2(n10781), .ZN(n10783) );
  AND2_X1 U13269 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12685) );
  INV_X1 U13270 ( .A(n12685), .ZN(n10782) );
  OAI211_X1 U13271 ( .C1(n15157), .C2(n10784), .A(n10783), .B(n10782), .ZN(
        n10785) );
  AOI21_X1 U13272 ( .B1(n11121), .B2(n13071), .A(n10785), .ZN(n10796) );
  NAND2_X1 U13273 ( .A1(n12985), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n10792) );
  INV_X1 U13274 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n10786) );
  MUX2_X1 U13275 ( .A(n10786), .B(P3_REG2_REG_12__SCAN_IN), .S(n12985), .Z(
        n10787) );
  INV_X1 U13276 ( .A(n10787), .ZN(n12989) );
  NAND2_X1 U13277 ( .A1(n10789), .A2(n10788), .ZN(n10791) );
  NAND2_X1 U13278 ( .A1(n10791), .A2(n10790), .ZN(n12990) );
  NAND2_X1 U13279 ( .A1(n12989), .A2(n12990), .ZN(n12988) );
  OAI21_X1 U13280 ( .B1(P3_REG2_REG_13__SCAN_IN), .B2(n10793), .A(n11116), 
        .ZN(n10794) );
  NAND2_X1 U13281 ( .A1(n10794), .A2(n15154), .ZN(n10795) );
  OAI211_X1 U13282 ( .C1(n10797), .C2(n13078), .A(n10796), .B(n10795), .ZN(
        P3_U3195) );
  NAND2_X1 U13283 ( .A1(n10800), .A2(SI_23_), .ZN(n11159) );
  OAI21_X1 U13284 ( .B1(SI_23_), .B2(n10800), .A(n11159), .ZN(n11156) );
  XNOR2_X1 U13285 ( .A(n11158), .B(n11156), .ZN(n11550) );
  INV_X1 U13286 ( .A(n11550), .ZN(n10802) );
  NAND2_X1 U13287 ( .A1(n14691), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n10801) );
  OAI211_X1 U13288 ( .C1(n10802), .C2(n14694), .A(n10801), .B(n12178), .ZN(
        P1_U3332) );
  INV_X1 U13289 ( .A(SI_25_), .ZN(n10806) );
  INV_X1 U13290 ( .A(n10803), .ZN(n10804) );
  OAI222_X1 U13291 ( .A1(n9579), .A2(n10806), .B1(P3_U3151), .B2(n10805), .C1(
        n12508), .C2(n10804), .ZN(P3_U3270) );
  INV_X1 U13292 ( .A(n10807), .ZN(n10808) );
  OAI222_X1 U13293 ( .A1(n9579), .A2(n10810), .B1(P3_U3151), .B2(n10809), .C1(
        n12508), .C2(n10808), .ZN(P3_U3269) );
  XNOR2_X1 U13294 ( .A(n10811), .B(n10812), .ZN(n15220) );
  NAND2_X1 U13295 ( .A1(n10814), .A2(n10813), .ZN(n10815) );
  NAND2_X1 U13296 ( .A1(n10815), .A2(n12932), .ZN(n10816) );
  NAND2_X1 U13297 ( .A1(n10817), .A2(n10816), .ZN(n10818) );
  NAND2_X1 U13298 ( .A1(n10818), .A2(n14762), .ZN(n10820) );
  AOI22_X1 U13299 ( .A1(n15192), .A2(n12972), .B1(n12970), .B2(n15195), .ZN(
        n10819) );
  OAI211_X1 U13300 ( .C1(n15177), .C2(n15220), .A(n10820), .B(n10819), .ZN(
        n15221) );
  MUX2_X1 U13301 ( .A(n15221), .B(P3_REG2_REG_8__SCAN_IN), .S(n15206), .Z(
        n10821) );
  INV_X1 U13302 ( .A(n10821), .ZN(n10825) );
  NOR2_X1 U13303 ( .A1(n10822), .A2(n15226), .ZN(n15222) );
  AOI22_X1 U13304 ( .A1(n14770), .A2(n15222), .B1(n15201), .B2(n10823), .ZN(
        n10824) );
  OAI211_X1 U13305 ( .C1(n15220), .C2(n13116), .A(n10825), .B(n10824), .ZN(
        P3_U3225) );
  NAND2_X1 U13306 ( .A1(n11550), .A2(n14078), .ZN(n10827) );
  NOR2_X1 U13307 ( .A1(n10826), .A2(P2_U3088), .ZN(n12491) );
  INV_X1 U13308 ( .A(n12491), .ZN(n12497) );
  OAI211_X1 U13309 ( .C1(n11551), .C2(n14086), .A(n10827), .B(n12497), .ZN(
        P2_U3304) );
  AND2_X1 U13310 ( .A1(n14828), .A2(n14256), .ZN(n10828) );
  NAND2_X1 U13311 ( .A1(n10830), .A2(n11913), .ZN(n10833) );
  AOI22_X1 U13312 ( .A1(n12116), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n11366), 
        .B2(n10831), .ZN(n10832) );
  XNOR2_X1 U13313 ( .A(n14734), .B(n14255), .ZN(n12145) );
  NAND2_X1 U13314 ( .A1(n14721), .A2(n14726), .ZN(n10835) );
  OR2_X1 U13315 ( .A1(n14734), .A2(n14255), .ZN(n10834) );
  NAND2_X1 U13316 ( .A1(n10835), .A2(n10834), .ZN(n10967) );
  NAND2_X1 U13317 ( .A1(n10836), .A2(n11913), .ZN(n10839) );
  AOI22_X1 U13318 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n12116), .B1(n10837), 
        .B2(n11366), .ZN(n10838) );
  NAND2_X1 U13319 ( .A1(n8996), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n10847) );
  OR2_X1 U13320 ( .A1(n9229), .A2(n10855), .ZN(n10846) );
  NAND2_X1 U13321 ( .A1(n10841), .A2(n10840), .ZN(n10842) );
  NAND2_X1 U13322 ( .A1(n10857), .A2(n10842), .ZN(n11217) );
  OR2_X1 U13323 ( .A1(n6575), .A2(n11217), .ZN(n10845) );
  OR2_X1 U13324 ( .A1(n11919), .A2(n10843), .ZN(n10844) );
  NAND4_X1 U13325 ( .A1(n10847), .A2(n10846), .A3(n10845), .A4(n10844), .ZN(
        n14254) );
  XNOR2_X1 U13326 ( .A(n14835), .B(n11212), .ZN(n12144) );
  XNOR2_X1 U13327 ( .A(n10967), .B(n12144), .ZN(n14840) );
  AOI21_X1 U13328 ( .B1(n14735), .B2(n14835), .A(n14924), .ZN(n10848) );
  OR2_X2 U13329 ( .A1(n14835), .A2(n14735), .ZN(n10976) );
  NAND2_X1 U13330 ( .A1(n10848), .A2(n10976), .ZN(n14836) );
  NOR2_X1 U13331 ( .A1(n14828), .A2(n14808), .ZN(n10850) );
  OR2_X1 U13332 ( .A1(n14734), .A2(n14819), .ZN(n10852) );
  NAND2_X1 U13333 ( .A1(n14722), .A2(n10852), .ZN(n10854) );
  INV_X1 U13334 ( .A(n12144), .ZN(n10853) );
  OR2_X1 U13335 ( .A1(n10854), .A2(n10853), .ZN(n14833) );
  NAND2_X1 U13336 ( .A1(n10854), .A2(n10853), .ZN(n10974) );
  NAND3_X1 U13337 ( .A1(n14833), .A2(n14480), .A3(n10974), .ZN(n10869) );
  NOR2_X1 U13338 ( .A1(n14544), .A2(n10855), .ZN(n10867) );
  NAND2_X1 U13339 ( .A1(n11381), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n10863) );
  OR2_X1 U13340 ( .A1(n9229), .A2(n10856), .ZN(n10862) );
  NAND2_X1 U13341 ( .A1(n10857), .A2(n14112), .ZN(n10858) );
  NAND2_X1 U13342 ( .A1(n10979), .A2(n10858), .ZN(n14117) );
  OR2_X1 U13343 ( .A1(n14117), .A2(n6575), .ZN(n10861) );
  OR2_X1 U13344 ( .A1(n11919), .A2(n10859), .ZN(n10860) );
  NAND2_X1 U13345 ( .A1(n14255), .A2(n14394), .ZN(n10864) );
  OAI21_X1 U13346 ( .B1(n11780), .B2(n14637), .A(n10864), .ZN(n14834) );
  INV_X1 U13347 ( .A(n14834), .ZN(n10865) );
  OAI22_X1 U13348 ( .A1(n14743), .A2(n10865), .B1(n11217), .B2(n14541), .ZN(
        n10866) );
  AOI211_X1 U13349 ( .C1(n14835), .C2(n14733), .A(n10867), .B(n10866), .ZN(
        n10868) );
  OAI211_X1 U13350 ( .C1(n14836), .C2(n14486), .A(n10869), .B(n10868), .ZN(
        n10870) );
  AOI21_X1 U13351 ( .B1(n14474), .B2(n14840), .A(n10870), .ZN(n10871) );
  INV_X1 U13352 ( .A(n10871), .ZN(P1_U3280) );
  AOI211_X1 U13353 ( .C1(n10874), .C2(n14012), .A(n10873), .B(n10872), .ZN(
        n10877) );
  AOI22_X1 U13354 ( .A1(n6593), .A2(n13992), .B1(P2_REG1_REG_14__SCAN_IN), 
        .B2(n15109), .ZN(n10875) );
  OAI21_X1 U13355 ( .B1(n10877), .B2(n15109), .A(n10875), .ZN(P2_U3513) );
  AOI22_X1 U13356 ( .A1(n6593), .A2(n14051), .B1(P2_REG0_REG_14__SCAN_IN), 
        .B2(n15104), .ZN(n10876) );
  OAI21_X1 U13357 ( .B1(n10877), .B2(n15104), .A(n10876), .ZN(P2_U3472) );
  NAND2_X1 U13358 ( .A1(n10878), .A2(n10886), .ZN(n10879) );
  NAND2_X1 U13359 ( .A1(n10880), .A2(n10879), .ZN(n15229) );
  NAND2_X1 U13360 ( .A1(n10881), .A2(n10992), .ZN(n10991) );
  NAND2_X1 U13361 ( .A1(n10991), .A2(n10882), .ZN(n10887) );
  AND2_X1 U13362 ( .A1(n10884), .A2(n10883), .ZN(n10885) );
  OAI211_X1 U13363 ( .C1(n10887), .C2(n10886), .A(n10885), .B(n14762), .ZN(
        n10889) );
  AOI22_X1 U13364 ( .A1(n15195), .A2(n12968), .B1(n12970), .B2(n15192), .ZN(
        n10888) );
  OAI211_X1 U13365 ( .C1(n15177), .C2(n15229), .A(n10889), .B(n10888), .ZN(
        n15231) );
  NAND2_X1 U13366 ( .A1(n15231), .A2(n15204), .ZN(n10893) );
  INV_X1 U13367 ( .A(n12597), .ZN(n10890) );
  OAI22_X1 U13368 ( .A1(n15204), .A2(n10339), .B1(n10890), .B2(n15169), .ZN(
        n10891) );
  AOI21_X1 U13369 ( .B1(n11101), .B2(n12588), .A(n10891), .ZN(n10892) );
  OAI211_X1 U13370 ( .C1(n15229), .C2(n13116), .A(n10893), .B(n10892), .ZN(
        P3_U3223) );
  XNOR2_X1 U13371 ( .A(n11256), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n10895) );
  NOR2_X1 U13372 ( .A1(n10896), .A2(n10895), .ZN(n11255) );
  AOI211_X1 U13373 ( .C1(n10896), .C2(n10895), .A(n15046), .B(n11255), .ZN(
        n10910) );
  INV_X1 U13374 ( .A(n10899), .ZN(n10904) );
  NAND2_X1 U13375 ( .A1(n10908), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n10897) );
  OAI211_X1 U13376 ( .C1(P2_REG2_REG_17__SCAN_IN), .C2(n10908), .A(n10898), 
        .B(n10897), .ZN(n10903) );
  NAND2_X1 U13377 ( .A1(n10899), .A2(n10898), .ZN(n10902) );
  NAND2_X1 U13378 ( .A1(n11256), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11250) );
  OAI21_X1 U13379 ( .B1(n11256), .B2(P2_REG2_REG_17__SCAN_IN), .A(n11250), 
        .ZN(n10900) );
  INV_X1 U13380 ( .A(n10900), .ZN(n10901) );
  NAND2_X1 U13381 ( .A1(n10902), .A2(n10901), .ZN(n11251) );
  OAI211_X1 U13382 ( .C1(n10904), .C2(n10903), .A(n11251), .B(n15039), .ZN(
        n10907) );
  AND2_X1 U13383 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n10905) );
  AOI21_X1 U13384 ( .B1(n14987), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n10905), 
        .ZN(n10906) );
  OAI211_X1 U13385 ( .C1(n14993), .C2(n10908), .A(n10907), .B(n10906), .ZN(
        n10909) );
  OR2_X1 U13386 ( .A1(n10910), .A2(n10909), .ZN(P2_U3231) );
  AOI211_X1 U13387 ( .C1(n14012), .C2(n10913), .A(n10912), .B(n10911), .ZN(
        n10916) );
  MUX2_X1 U13388 ( .A(n10914), .B(n10916), .S(n15112), .Z(n10915) );
  OAI21_X1 U13389 ( .B1(n10919), .B2(n14015), .A(n10915), .ZN(P2_U3514) );
  MUX2_X1 U13390 ( .A(n10917), .B(n10916), .S(n15106), .Z(n10918) );
  OAI21_X1 U13391 ( .B1(n10919), .B2(n14064), .A(n10918), .ZN(P2_U3475) );
  OR2_X1 U13392 ( .A1(n12300), .A2(n13547), .ZN(n10922) );
  NAND2_X1 U13393 ( .A1(n11168), .A2(n12393), .ZN(n10925) );
  AOI22_X1 U13394 ( .A1(n11505), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n10923), 
        .B2(n11504), .ZN(n10924) );
  INV_X1 U13395 ( .A(n13546), .ZN(n12310) );
  XNOR2_X1 U13396 ( .A(n12308), .B(n12310), .ZN(n12471) );
  NAND2_X1 U13397 ( .A1(n10926), .A2(n7225), .ZN(n10927) );
  NAND2_X1 U13398 ( .A1(n11145), .A2(n10927), .ZN(n11201) );
  OR2_X2 U13399 ( .A1(n10928), .A2(n12470), .ZN(n10931) );
  NAND2_X1 U13400 ( .A1(n12300), .A2(n10929), .ZN(n10930) );
  AOI21_X1 U13401 ( .B1(n10932), .B2(n12471), .A(n13875), .ZN(n10933) );
  NAND2_X1 U13402 ( .A1(n10933), .A2(n11142), .ZN(n11200) );
  NAND2_X1 U13403 ( .A1(n10934), .A2(n11084), .ZN(n10935) );
  AND2_X1 U13404 ( .A1(n11075), .A2(n10935), .ZN(n11150) );
  NAND2_X1 U13405 ( .A1(n11150), .A2(n6638), .ZN(n10940) );
  INV_X1 U13406 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14013) );
  NAND2_X1 U13407 ( .A1(n11619), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n10937) );
  NAND2_X1 U13408 ( .A1(n11618), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n10936) );
  OAI211_X1 U13409 ( .C1(n14013), .C2(n11609), .A(n10937), .B(n10936), .ZN(
        n10938) );
  INV_X1 U13410 ( .A(n10938), .ZN(n10939) );
  NAND2_X1 U13411 ( .A1(n10940), .A2(n10939), .ZN(n13545) );
  AND2_X1 U13412 ( .A1(n13547), .A2(n13518), .ZN(n10941) );
  AOI21_X1 U13413 ( .B1(n13545), .B2(n13517), .A(n10941), .ZN(n11197) );
  OAI211_X1 U13414 ( .C1(n13825), .C2(n11108), .A(n11200), .B(n11197), .ZN(
        n10942) );
  NAND2_X1 U13415 ( .A1(n10942), .A2(n13868), .ZN(n10950) );
  INV_X1 U13416 ( .A(n12308), .ZN(n10946) );
  OAI21_X1 U13417 ( .B1(n10946), .B2(n10943), .A(n9326), .ZN(n10944) );
  OR2_X1 U13418 ( .A1(n11147), .A2(n10944), .ZN(n11198) );
  INV_X1 U13419 ( .A(n11198), .ZN(n10948) );
  INV_X1 U13420 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n10945) );
  OAI22_X1 U13421 ( .A1(n10946), .A2(n15069), .B1(n10945), .B2(n13868), .ZN(
        n10947) );
  AOI21_X1 U13422 ( .B1(n10948), .B2(n15064), .A(n10947), .ZN(n10949) );
  OAI211_X1 U13423 ( .C1(n11201), .C2(n13871), .A(n10950), .B(n10949), .ZN(
        P2_U3249) );
  XNOR2_X1 U13424 ( .A(n12614), .B(n15164), .ZN(n12512) );
  XNOR2_X1 U13425 ( .A(n12512), .B(n12970), .ZN(n10959) );
  INV_X1 U13426 ( .A(n10951), .ZN(n10952) );
  NAND2_X1 U13427 ( .A1(n10952), .A2(n12971), .ZN(n10953) );
  INV_X1 U13428 ( .A(n10958), .ZN(n10956) );
  INV_X1 U13429 ( .A(n12514), .ZN(n10957) );
  AOI21_X1 U13430 ( .B1(n10959), .B2(n10958), .A(n10957), .ZN(n10966) );
  OAI22_X1 U13431 ( .A1(n12720), .A2(n15164), .B1(n10960), .B2(n12719), .ZN(
        n10961) );
  AOI211_X1 U13432 ( .C1(n12717), .C2(n12969), .A(n10962), .B(n10961), .ZN(
        n10965) );
  NAND2_X1 U13433 ( .A1(n12729), .A2(n10963), .ZN(n10964) );
  OAI211_X1 U13434 ( .C1(n10966), .C2(n12739), .A(n10965), .B(n10964), .ZN(
        P3_U3171) );
  NAND2_X1 U13435 ( .A1(n10968), .A2(n11913), .ZN(n10971) );
  AOI22_X1 U13436 ( .A1(n10969), .A2(n11366), .B1(P2_DATAO_REG_14__SCAN_IN), 
        .B2(n12116), .ZN(n10970) );
  NAND2_X1 U13437 ( .A1(n14119), .A2(n11780), .ZN(n12022) );
  OAI21_X1 U13438 ( .B1(n7421), .B2(n10972), .A(n11177), .ZN(n11041) );
  OR2_X1 U13439 ( .A1(n14835), .A2(n11212), .ZN(n10973) );
  XOR2_X1 U13440 ( .A(n12147), .B(n11184), .Z(n11043) );
  NAND2_X1 U13441 ( .A1(n11043), .A2(n14480), .ZN(n10990) );
  NAND2_X1 U13442 ( .A1(n14119), .A2(n10976), .ZN(n10975) );
  NAND2_X1 U13443 ( .A1(n10975), .A2(n14736), .ZN(n10977) );
  OR2_X1 U13444 ( .A1(n10977), .A2(n14531), .ZN(n11039) );
  INV_X1 U13445 ( .A(n11039), .ZN(n10988) );
  INV_X1 U13446 ( .A(n14119), .ZN(n11779) );
  INV_X1 U13447 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n10978) );
  AND2_X1 U13448 ( .A1(n10979), .A2(n10978), .ZN(n10980) );
  OR2_X1 U13449 ( .A1(n10980), .A2(n11172), .ZN(n14542) );
  OAI22_X1 U13450 ( .A1(n14542), .A2(n6575), .B1(n11919), .B2(n14898), .ZN(
        n10981) );
  INV_X1 U13451 ( .A(n10981), .ZN(n10983) );
  AOI22_X1 U13452 ( .A1(n11459), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n11381), 
        .B2(P1_REG0_REG_15__SCAN_IN), .ZN(n10982) );
  OAI22_X1 U13453 ( .A1(n14113), .A2(n14637), .B1(n11212), .B2(n14517), .ZN(
        n11038) );
  INV_X1 U13454 ( .A(n11038), .ZN(n10984) );
  OAI22_X1 U13455 ( .A1(n14743), .A2(n10984), .B1(n14117), .B2(n14541), .ZN(
        n10985) );
  AOI21_X1 U13456 ( .B1(n14743), .B2(P1_REG2_REG_14__SCAN_IN), .A(n10985), 
        .ZN(n10986) );
  OAI21_X1 U13457 ( .B1(n11779), .B2(n14506), .A(n10986), .ZN(n10987) );
  AOI21_X1 U13458 ( .B1(n10988), .B2(n14739), .A(n10987), .ZN(n10989) );
  OAI211_X1 U13459 ( .C1(n11041), .C2(n14546), .A(n10990), .B(n10989), .ZN(
        P1_U3279) );
  OAI211_X1 U13460 ( .C1(n10881), .C2(n10992), .A(n10991), .B(n14762), .ZN(
        n10994) );
  AOI22_X1 U13461 ( .A1(n15192), .A2(n12971), .B1(n12969), .B2(n15195), .ZN(
        n10993) );
  AND2_X1 U13462 ( .A1(n10994), .A2(n10993), .ZN(n15160) );
  XNOR2_X1 U13463 ( .A(n10995), .B(n12936), .ZN(n15159) );
  NAND2_X1 U13464 ( .A1(n15159), .A2(n14798), .ZN(n10996) );
  AND2_X1 U13465 ( .A1(n15160), .A2(n10996), .ZN(n10999) );
  INV_X1 U13466 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n10997) );
  MUX2_X1 U13467 ( .A(n10999), .B(n10997), .S(n15234), .Z(n10998) );
  OAI21_X1 U13468 ( .B1(n13384), .B2(n15164), .A(n10998), .ZN(P3_U3417) );
  INV_X1 U13469 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11000) );
  MUX2_X1 U13470 ( .A(n11000), .B(n10999), .S(n15240), .Z(n11001) );
  OAI21_X1 U13471 ( .B1(n13334), .B2(n15164), .A(n11001), .ZN(P3_U3468) );
  INV_X1 U13472 ( .A(n11002), .ZN(n11004) );
  NOR2_X1 U13473 ( .A1(n14807), .A2(n11879), .ZN(n11006) );
  AOI21_X1 U13474 ( .B1(n14962), .B2(n11825), .A(n11006), .ZN(n11010) );
  AOI22_X1 U13475 ( .A1(n14962), .A2(n11870), .B1(n11825), .B2(n14258), .ZN(
        n11007) );
  XNOR2_X1 U13476 ( .A(n11007), .B(n11881), .ZN(n14874) );
  INV_X1 U13477 ( .A(n11008), .ZN(n11009) );
  NAND2_X1 U13478 ( .A1(n14806), .A2(n11870), .ZN(n11012) );
  NAND2_X1 U13479 ( .A1(n14257), .A2(n6423), .ZN(n11011) );
  NAND2_X1 U13480 ( .A1(n11012), .A2(n11011), .ZN(n11013) );
  XNOR2_X1 U13481 ( .A(n11013), .B(n11881), .ZN(n11021) );
  NOR2_X1 U13482 ( .A1(n14872), .A2(n11879), .ZN(n11014) );
  AOI21_X1 U13483 ( .B1(n14806), .B2(n11825), .A(n11014), .ZN(n11019) );
  XNOR2_X1 U13484 ( .A(n11021), .B(n11019), .ZN(n14810) );
  NAND2_X1 U13485 ( .A1(n14828), .A2(n11870), .ZN(n11016) );
  NAND2_X1 U13486 ( .A1(n14256), .A2(n6423), .ZN(n11015) );
  NAND2_X1 U13487 ( .A1(n11016), .A2(n11015), .ZN(n11017) );
  XNOR2_X1 U13488 ( .A(n11017), .B(n11881), .ZN(n11025) );
  NOR2_X1 U13489 ( .A1(n14808), .A2(n11879), .ZN(n11018) );
  AOI21_X1 U13490 ( .B1(n14828), .B2(n11825), .A(n11018), .ZN(n11023) );
  XNOR2_X1 U13491 ( .A(n11025), .B(n11023), .ZN(n14820) );
  INV_X1 U13492 ( .A(n11019), .ZN(n11020) );
  NAND2_X1 U13493 ( .A1(n11021), .A2(n11020), .ZN(n14821) );
  INV_X1 U13494 ( .A(n11023), .ZN(n11024) );
  NOR2_X1 U13495 ( .A1(n14819), .A2(n11879), .ZN(n11027) );
  AOI21_X1 U13496 ( .B1(n14734), .B2(n11825), .A(n11027), .ZN(n11210) );
  NAND2_X1 U13497 ( .A1(n14734), .A2(n11870), .ZN(n11029) );
  NAND2_X1 U13498 ( .A1(n14255), .A2(n11825), .ZN(n11028) );
  NAND2_X1 U13499 ( .A1(n11029), .A2(n11028), .ZN(n11030) );
  XNOR2_X1 U13500 ( .A(n11030), .B(n11881), .ZN(n11207) );
  XOR2_X1 U13501 ( .A(n11210), .B(n11207), .Z(n11032) );
  AOI21_X1 U13502 ( .B1(n11031), .B2(n11032), .A(n14875), .ZN(n11033) );
  NAND2_X1 U13503 ( .A1(n11033), .A2(n11208), .ZN(n11037) );
  INV_X1 U13504 ( .A(n14233), .ZN(n14225) );
  OAI22_X1 U13505 ( .A1(n14808), .A2(n14517), .B1(n11212), .B2(n14637), .ZN(
        n14728) );
  NOR2_X1 U13506 ( .A1(n14883), .A2(n14730), .ZN(n11034) );
  AOI211_X1 U13507 ( .C1(n14225), .C2(n14728), .A(n11035), .B(n11034), .ZN(
        n11036) );
  OAI211_X1 U13508 ( .C1(n14745), .C2(n14239), .A(n11037), .B(n11036), .ZN(
        P1_U3224) );
  AOI21_X1 U13509 ( .B1(n14119), .B2(n14961), .A(n11038), .ZN(n11040) );
  OAI211_X1 U13510 ( .C1(n11041), .C2(n14969), .A(n11040), .B(n11039), .ZN(
        n11042) );
  AOI21_X1 U13511 ( .B1(n14832), .B2(n11043), .A(n11042), .ZN(n11046) );
  NAND2_X1 U13512 ( .A1(n14984), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11044) );
  OAI21_X1 U13513 ( .B1(n11046), .B2(n14984), .A(n11044), .ZN(P1_U3542) );
  NAND2_X1 U13514 ( .A1(n14975), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11045) );
  OAI21_X1 U13515 ( .B1(n11046), .B2(n14975), .A(n11045), .ZN(P1_U3501) );
  INV_X1 U13516 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n11047) );
  XNOR2_X1 U13517 ( .A(n14295), .B(n11047), .ZN(n14298) );
  INV_X1 U13518 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11050) );
  INV_X1 U13519 ( .A(n11048), .ZN(n11049) );
  OAI21_X1 U13520 ( .B1(n11054), .B2(n11050), .A(n11049), .ZN(n14297) );
  NAND2_X1 U13521 ( .A1(n14298), .A2(n14297), .ZN(n14296) );
  NAND2_X1 U13522 ( .A1(n14295), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n11051) );
  XNOR2_X1 U13523 ( .A(n14308), .B(n14307), .ZN(n11052) );
  INV_X1 U13524 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n11362) );
  NOR2_X1 U13525 ( .A1(n11362), .A2(n11052), .ZN(n14309) );
  AOI211_X1 U13526 ( .C1(n11052), .C2(n11362), .A(n14309), .B(n14323), .ZN(
        n11062) );
  INV_X1 U13527 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11056) );
  OAI21_X1 U13528 ( .B1(n11054), .B2(n10483), .A(n11053), .ZN(n14303) );
  NAND2_X1 U13529 ( .A1(n14300), .A2(n11056), .ZN(n11055) );
  OAI211_X1 U13530 ( .C1(n14300), .C2(n11056), .A(n14303), .B(n11055), .ZN(
        n14301) );
  OAI21_X1 U13531 ( .B1(n11056), .B2(n14300), .A(n14301), .ZN(n14313) );
  XNOR2_X1 U13532 ( .A(n14313), .B(n14307), .ZN(n11057) );
  NAND2_X1 U13533 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n11057), .ZN(n14316) );
  OAI211_X1 U13534 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n11057), .A(n14318), 
        .B(n14316), .ZN(n11060) );
  NAND2_X1 U13535 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14215)
         );
  INV_X1 U13536 ( .A(n14215), .ZN(n11058) );
  AOI21_X1 U13537 ( .B1(n14891), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n11058), 
        .ZN(n11059) );
  OAI211_X1 U13538 ( .C1(n14320), .C2(n14307), .A(n11060), .B(n11059), .ZN(
        n11061) );
  OR2_X1 U13539 ( .A1(n11062), .A2(n11061), .ZN(P1_U3261) );
  INV_X1 U13540 ( .A(n11063), .ZN(n11065) );
  XNOR2_X1 U13541 ( .A(n12308), .B(n13424), .ZN(n11088) );
  NAND2_X1 U13542 ( .A1(n13546), .A2(n13845), .ZN(n11068) );
  XNOR2_X1 U13543 ( .A(n11088), .B(n11068), .ZN(n11107) );
  NAND2_X1 U13544 ( .A1(n11088), .A2(n11068), .ZN(n11069) );
  NAND2_X1 U13545 ( .A1(n11353), .A2(n12393), .ZN(n11071) );
  AOI22_X1 U13546 ( .A1(n11505), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n11504), 
        .B2(n11256), .ZN(n11070) );
  XNOR2_X1 U13547 ( .A(n12314), .B(n6627), .ZN(n11671) );
  NAND2_X1 U13548 ( .A1(n13545), .A2(n13845), .ZN(n11672) );
  XNOR2_X1 U13549 ( .A(n11671), .B(n11672), .ZN(n11087) );
  INV_X1 U13550 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n11074) );
  NAND2_X1 U13551 ( .A1(n11075), .A2(n11074), .ZN(n11076) );
  NAND2_X1 U13552 ( .A1(n11233), .A2(n11076), .ZN(n13499) );
  OR2_X1 U13553 ( .A1(n13499), .A2(n11606), .ZN(n11082) );
  INV_X1 U13554 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n11079) );
  NAND2_X1 U13555 ( .A1(n11619), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n11078) );
  NAND2_X1 U13556 ( .A1(n11618), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n11077) );
  OAI211_X1 U13557 ( .C1(n11079), .C2(n11609), .A(n11078), .B(n11077), .ZN(
        n11080) );
  INV_X1 U13558 ( .A(n11080), .ZN(n11081) );
  NAND2_X1 U13559 ( .A1(n11082), .A2(n11081), .ZN(n13544) );
  AND2_X1 U13560 ( .A1(n13546), .A2(n13518), .ZN(n11083) );
  AOI21_X1 U13561 ( .B1(n13544), .B2(n13517), .A(n11083), .ZN(n11143) );
  OAI22_X1 U13562 ( .A1(n13503), .A2(n11143), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11084), .ZN(n11086) );
  NOR2_X1 U13563 ( .A1(n14065), .A2(n13525), .ZN(n11085) );
  AOI211_X1 U13564 ( .C1(n13522), .C2(n11150), .A(n11086), .B(n11085), .ZN(
        n11092) );
  INV_X1 U13565 ( .A(n11087), .ZN(n11090) );
  OAI22_X1 U13566 ( .A1(n11088), .A2(n13478), .B1(n12310), .B2(n13512), .ZN(
        n11089) );
  NAND3_X1 U13567 ( .A1(n11104), .A2(n11090), .A3(n11089), .ZN(n11091) );
  OAI211_X1 U13568 ( .C1(n11675), .C2(n13478), .A(n11092), .B(n11091), .ZN(
        P2_U3200) );
  XNOR2_X1 U13569 ( .A(n11093), .B(n11096), .ZN(n14791) );
  NAND2_X1 U13570 ( .A1(n11095), .A2(n11094), .ZN(n11097) );
  XNOR2_X1 U13571 ( .A(n11097), .B(n11096), .ZN(n11098) );
  OAI222_X1 U13572 ( .A1(n14776), .A2(n6878), .B1(n14778), .B2(n12700), .C1(
        n11098), .C2(n15198), .ZN(n14793) );
  NAND2_X1 U13573 ( .A1(n14793), .A2(n15204), .ZN(n11103) );
  INV_X1 U13574 ( .A(n12637), .ZN(n11099) );
  OAI22_X1 U13575 ( .A1(n15204), .A2(n10786), .B1(n11099), .B2(n15169), .ZN(
        n11100) );
  AOI21_X1 U13576 ( .B1(n11101), .B2(n12634), .A(n11100), .ZN(n11102) );
  OAI211_X1 U13577 ( .C1(n13207), .C2(n14791), .A(n11103), .B(n11102), .ZN(
        P3_U3221) );
  INV_X1 U13578 ( .A(n11104), .ZN(n11105) );
  AOI21_X1 U13579 ( .B1(n11107), .B2(n11106), .A(n11105), .ZN(n11113) );
  NOR2_X1 U13580 ( .A1(n13495), .A2(n11108), .ZN(n11111) );
  OAI22_X1 U13581 ( .A1(n13503), .A2(n11197), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11109), .ZN(n11110) );
  AOI211_X1 U13582 ( .C1(n12308), .C2(n13510), .A(n11111), .B(n11110), .ZN(
        n11112) );
  OAI21_X1 U13583 ( .B1(n11113), .B2(n13478), .A(n11112), .ZN(P2_U3198) );
  INV_X1 U13584 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13740) );
  OR2_X1 U13585 ( .A1(n11122), .A2(n13740), .ZN(n11278) );
  NAND2_X1 U13586 ( .A1(n11122), .A2(n13740), .ZN(n11114) );
  AND2_X1 U13587 ( .A1(n11278), .A2(n11114), .ZN(n11267) );
  NAND2_X1 U13588 ( .A1(n11127), .A2(n11115), .ZN(n11117) );
  XOR2_X1 U13589 ( .A(n11267), .B(n11266), .Z(n11140) );
  INV_X1 U13590 ( .A(n11118), .ZN(n11120) );
  INV_X1 U13591 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13332) );
  OR2_X1 U13592 ( .A1(n11122), .A2(n13332), .ZN(n11277) );
  NAND2_X1 U13593 ( .A1(n11122), .A2(n13332), .ZN(n11123) );
  AND2_X1 U13594 ( .A1(n11277), .A2(n11123), .ZN(n11131) );
  MUX2_X1 U13595 ( .A(n11267), .B(n11131), .S(n13037), .Z(n11124) );
  NAND2_X1 U13596 ( .A1(n11125), .A2(n11124), .ZN(n11280) );
  INV_X1 U13597 ( .A(n13078), .ZN(n15146) );
  OAI211_X1 U13598 ( .C1(n11125), .C2(n11124), .A(n11280), .B(n15146), .ZN(
        n11138) );
  NAND2_X1 U13599 ( .A1(n11127), .A2(n11126), .ZN(n11129) );
  NAND2_X1 U13600 ( .A1(n11129), .A2(n11128), .ZN(n11130) );
  NAND2_X1 U13601 ( .A1(n11130), .A2(n11131), .ZN(n11271) );
  OAI21_X1 U13602 ( .B1(n11131), .B2(n11130), .A(n11271), .ZN(n11136) );
  INV_X1 U13603 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n11132) );
  NOR2_X1 U13604 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11132), .ZN(n12575) );
  AOI21_X1 U13605 ( .B1(n15113), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12575), 
        .ZN(n11133) );
  OAI21_X1 U13606 ( .B1(n15150), .B2(n11134), .A(n11133), .ZN(n11135) );
  AOI21_X1 U13607 ( .B1(n11136), .B2(n13023), .A(n11135), .ZN(n11137) );
  OAI211_X1 U13608 ( .C1(n11140), .C2(n11139), .A(n11138), .B(n11137), .ZN(
        P3_U3196) );
  INV_X1 U13609 ( .A(n13545), .ZN(n11230) );
  XNOR2_X1 U13610 ( .A(n12314), .B(n11230), .ZN(n12473) );
  OR2_X1 U13611 ( .A1(n12308), .A2(n12310), .ZN(n11141) );
  XOR2_X1 U13612 ( .A(n12473), .B(n11229), .Z(n11144) );
  OAI21_X1 U13613 ( .B1(n11144), .B2(n13875), .A(n11143), .ZN(n14009) );
  INV_X1 U13614 ( .A(n14009), .ZN(n11155) );
  INV_X1 U13615 ( .A(n12473), .ZN(n11146) );
  XNOR2_X1 U13616 ( .A(n11222), .B(n11146), .ZN(n14011) );
  INV_X1 U13617 ( .A(n11147), .ZN(n11149) );
  INV_X1 U13618 ( .A(n11242), .ZN(n11148) );
  AOI211_X1 U13619 ( .C1(n12314), .C2(n11149), .A(n6649), .B(n11148), .ZN(
        n14010) );
  NAND2_X1 U13620 ( .A1(n14010), .A2(n15064), .ZN(n11152) );
  AOI22_X1 U13621 ( .A1(n15075), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n11150), 
        .B2(n15062), .ZN(n11151) );
  OAI211_X1 U13622 ( .C1(n14065), .C2(n15069), .A(n11152), .B(n11151), .ZN(
        n11153) );
  AOI21_X1 U13623 ( .B1(n15072), .B2(n14011), .A(n11153), .ZN(n11154) );
  OAI21_X1 U13624 ( .B1(n11155), .B2(n15075), .A(n11154), .ZN(P2_U3248) );
  INV_X1 U13625 ( .A(n11156), .ZN(n11157) );
  MUX2_X1 U13626 ( .A(n11163), .B(n11565), .S(n11907), .Z(n11160) );
  NAND2_X1 U13627 ( .A1(n11161), .A2(n11160), .ZN(n11162) );
  INV_X1 U13628 ( .A(n11564), .ZN(n11166) );
  OAI222_X1 U13629 ( .A1(n11164), .A2(P1_U3086), .B1(n14694), .B2(n11166), 
        .C1(n11163), .C2(n14684), .ZN(P1_U3331) );
  INV_X1 U13630 ( .A(n11165), .ZN(n11167) );
  OAI222_X1 U13631 ( .A1(P2_U3088), .A2(n11167), .B1(n14086), .B2(n11565), 
        .C1(n14088), .C2(n11166), .ZN(P2_U3303) );
  NAND2_X1 U13632 ( .A1(n11168), .A2(n11913), .ZN(n11171) );
  AOI22_X1 U13633 ( .A1(n12116), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11366), 
        .B2(n11169), .ZN(n11170) );
  NOR2_X1 U13634 ( .A1(n11172), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11173) );
  OR2_X1 U13635 ( .A1(n11186), .A2(n11173), .ZN(n14171) );
  AOI22_X1 U13636 ( .A1(n11459), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n11381), 
        .B2(P1_REG0_REG_16__SCAN_IN), .ZN(n11175) );
  INV_X1 U13637 ( .A(n11919), .ZN(n11320) );
  NAND2_X1 U13638 ( .A1(n11320), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11174) );
  OAI211_X1 U13639 ( .C1(n14171), .C2(n6575), .A(n11175), .B(n11174), .ZN(
        n14251) );
  INV_X1 U13640 ( .A(n14251), .ZN(n14518) );
  XNOR2_X1 U13641 ( .A(n14173), .B(n14518), .ZN(n12149) );
  INV_X1 U13642 ( .A(n11780), .ZN(n14253) );
  NAND2_X1 U13643 ( .A1(n14119), .A2(n14253), .ZN(n11176) );
  NAND2_X1 U13644 ( .A1(n11178), .A2(n11913), .ZN(n11180) );
  AOI22_X1 U13645 ( .A1(n12116), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11366), 
        .B2(n14902), .ZN(n11179) );
  NAND2_X1 U13646 ( .A1(n14653), .A2(n14113), .ZN(n12023) );
  INV_X1 U13647 ( .A(n14534), .ZN(n11181) );
  INV_X1 U13648 ( .A(n14113), .ZN(n14252) );
  OR2_X1 U13649 ( .A1(n14653), .A2(n14252), .ZN(n11182) );
  XOR2_X1 U13650 ( .A(n11351), .B(n12149), .Z(n14651) );
  INV_X1 U13651 ( .A(n12149), .ZN(n11185) );
  OAI21_X1 U13652 ( .B1(n6544), .B2(n11185), .A(n11444), .ZN(n14649) );
  INV_X1 U13653 ( .A(n14653), .ZN(n14240) );
  AND2_X1 U13654 ( .A1(n14531), .A2(n14240), .ZN(n14532) );
  NAND2_X1 U13655 ( .A1(n14532), .A2(n14647), .ZN(n14519) );
  OAI211_X1 U13656 ( .C1(n14532), .C2(n14647), .A(n14736), .B(n14519), .ZN(
        n14646) );
  NOR2_X1 U13657 ( .A1(n11186), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11187) );
  OR2_X1 U13658 ( .A1(n11360), .A2(n11187), .ZN(n14522) );
  AOI22_X1 U13659 ( .A1(n11459), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n11381), 
        .B2(P1_REG0_REG_17__SCAN_IN), .ZN(n11189) );
  NAND2_X1 U13660 ( .A1(n11320), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n11188) );
  OAI211_X1 U13661 ( .C1(n14522), .C2(n6575), .A(n11189), .B(n11188), .ZN(
        n14250) );
  NAND2_X1 U13662 ( .A1(n14250), .A2(n14921), .ZN(n11191) );
  OR2_X1 U13663 ( .A1(n14113), .A2(n14517), .ZN(n11190) );
  NAND2_X1 U13664 ( .A1(n11191), .A2(n11190), .ZN(n14169) );
  INV_X1 U13665 ( .A(n14169), .ZN(n14645) );
  OAI22_X1 U13666 ( .A1(n14743), .A2(n14645), .B1(n14171), .B2(n14541), .ZN(
        n11193) );
  NOR2_X1 U13667 ( .A1(n14647), .A2(n14506), .ZN(n11192) );
  AOI211_X1 U13668 ( .C1(n14743), .C2(P1_REG2_REG_16__SCAN_IN), .A(n11193), 
        .B(n11192), .ZN(n11194) );
  OAI21_X1 U13669 ( .B1(n14486), .B2(n14646), .A(n11194), .ZN(n11195) );
  AOI21_X1 U13670 ( .B1(n14649), .B2(n14480), .A(n11195), .ZN(n11196) );
  OAI21_X1 U13671 ( .B1(n14651), .B2(n14546), .A(n11196), .ZN(P1_U3277) );
  AND2_X1 U13672 ( .A1(n11198), .A2(n11197), .ZN(n11199) );
  OAI211_X1 U13673 ( .C1(n11201), .C2(n15093), .A(n11200), .B(n11199), .ZN(
        n11204) );
  MUX2_X1 U13674 ( .A(n11204), .B(P2_REG1_REG_16__SCAN_IN), .S(n15109), .Z(
        n11202) );
  AOI21_X1 U13675 ( .B1(n13992), .B2(n12308), .A(n11202), .ZN(n11203) );
  INV_X1 U13676 ( .A(n11203), .ZN(P2_U3515) );
  MUX2_X1 U13677 ( .A(n11204), .B(P2_REG0_REG_16__SCAN_IN), .S(n15104), .Z(
        n11205) );
  AOI21_X1 U13678 ( .B1(n14051), .B2(n12308), .A(n11205), .ZN(n11206) );
  INV_X1 U13679 ( .A(n11206), .ZN(P2_U3478) );
  INV_X1 U13680 ( .A(n14835), .ZN(n12017) );
  INV_X1 U13681 ( .A(n11207), .ZN(n11209) );
  OAI22_X1 U13682 ( .A1(n12017), .A2(n11880), .B1(n11212), .B2(n8975), .ZN(
        n11211) );
  XNOR2_X1 U13683 ( .A(n11211), .B(n11881), .ZN(n11784) );
  NOR2_X1 U13684 ( .A1(n11212), .A2(n11879), .ZN(n11213) );
  AOI21_X1 U13685 ( .B1(n14835), .B2(n6423), .A(n11213), .ZN(n11786) );
  XNOR2_X1 U13686 ( .A(n11784), .B(n11786), .ZN(n11214) );
  OAI211_X1 U13687 ( .C1(n11215), .C2(n11214), .A(n11785), .B(n14809), .ZN(
        n11221) );
  OAI21_X1 U13688 ( .B1(n14871), .B2(n11780), .A(n11216), .ZN(n11219) );
  NOR2_X1 U13689 ( .A1(n14883), .A2(n11217), .ZN(n11218) );
  AOI211_X1 U13690 ( .C1(n14115), .C2(n14255), .A(n11219), .B(n11218), .ZN(
        n11220) );
  OAI211_X1 U13691 ( .C1(n12017), .C2(n14239), .A(n11221), .B(n11220), .ZN(
        P1_U3234) );
  NAND2_X1 U13692 ( .A1(n11222), .A2(n12473), .ZN(n11224) );
  NAND2_X1 U13693 ( .A1(n12314), .A2(n13545), .ZN(n11223) );
  NAND2_X1 U13694 ( .A1(n11357), .A2(n12393), .ZN(n11227) );
  AOI22_X1 U13695 ( .A1(n11505), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n11504), 
        .B2(n11225), .ZN(n11226) );
  INV_X1 U13696 ( .A(n13544), .ZN(n13445) );
  XNOR2_X1 U13697 ( .A(n14006), .B(n13445), .ZN(n12475) );
  XNOR2_X1 U13698 ( .A(n11634), .B(n12475), .ZN(n14008) );
  NOR2_X1 U13699 ( .A1(n12314), .A2(n11230), .ZN(n11228) );
  INV_X1 U13700 ( .A(n12475), .ZN(n11633) );
  NAND2_X1 U13701 ( .A1(n11231), .A2(n11633), .ZN(n11502) );
  OAI211_X1 U13702 ( .C1(n11231), .C2(n11633), .A(n11502), .B(n13891), .ZN(
        n11241) );
  INV_X1 U13703 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n11232) );
  NAND2_X1 U13704 ( .A1(n11233), .A2(n11232), .ZN(n11234) );
  AND2_X1 U13705 ( .A1(n11516), .A2(n11234), .ZN(n13900) );
  NAND2_X1 U13706 ( .A1(n13900), .A2(n6638), .ZN(n11239) );
  INV_X1 U13707 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14002) );
  NAND2_X1 U13708 ( .A1(n11619), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n11236) );
  NAND2_X1 U13709 ( .A1(n11618), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n11235) );
  OAI211_X1 U13710 ( .C1(n14002), .C2(n11609), .A(n11236), .B(n11235), .ZN(
        n11237) );
  INV_X1 U13711 ( .A(n11237), .ZN(n11238) );
  NAND2_X1 U13712 ( .A1(n11239), .A2(n11238), .ZN(n13543) );
  AND2_X1 U13713 ( .A1(n13545), .A2(n13518), .ZN(n11240) );
  AOI21_X1 U13714 ( .B1(n13543), .B2(n13517), .A(n11240), .ZN(n13504) );
  NAND2_X1 U13715 ( .A1(n11241), .A2(n13504), .ZN(n14004) );
  AOI21_X1 U13716 ( .B1(n14006), .B2(n11242), .A(n6649), .ZN(n11243) );
  AND2_X1 U13717 ( .A1(n11243), .A2(n13898), .ZN(n14005) );
  NAND2_X1 U13718 ( .A1(n14005), .A2(n13923), .ZN(n11247) );
  NAND2_X1 U13719 ( .A1(n15075), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n11244) );
  OAI21_X1 U13720 ( .B1(n13825), .B2(n13499), .A(n11244), .ZN(n11245) );
  AOI21_X1 U13721 ( .B1(n14006), .B2(n13927), .A(n11245), .ZN(n11246) );
  NAND2_X1 U13722 ( .A1(n11247), .A2(n11246), .ZN(n11248) );
  AOI21_X1 U13723 ( .B1(n14004), .B2(n13868), .A(n11248), .ZN(n11249) );
  OAI21_X1 U13724 ( .B1(n14008), .B2(n13871), .A(n11249), .ZN(P2_U3247) );
  AND2_X1 U13725 ( .A1(n11253), .A2(n11261), .ZN(n13568) );
  INV_X1 U13726 ( .A(n13568), .ZN(n11252) );
  OAI21_X1 U13727 ( .B1(n11253), .B2(n11261), .A(n11252), .ZN(n11254) );
  AOI21_X1 U13728 ( .B1(n11254), .B2(P2_REG2_REG_18__SCAN_IN), .A(n13567), 
        .ZN(n11265) );
  NOR2_X1 U13729 ( .A1(n11257), .A2(n11261), .ZN(n13564) );
  AOI21_X1 U13730 ( .B1(n11257), .B2(n11261), .A(n13564), .ZN(n11259) );
  AND2_X1 U13731 ( .A1(n11259), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n13565) );
  INV_X1 U13732 ( .A(n13565), .ZN(n11258) );
  OAI211_X1 U13733 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n11259), .A(n11258), 
        .B(n15003), .ZN(n11264) );
  NAND2_X1 U13734 ( .A1(n14987), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n11260) );
  NAND2_X1 U13735 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13501)
         );
  OAI211_X1 U13736 ( .C1(n14993), .C2(n11261), .A(n11260), .B(n13501), .ZN(
        n11262) );
  INV_X1 U13737 ( .A(n11262), .ZN(n11263) );
  OAI211_X1 U13738 ( .C1(n11265), .C2(n15054), .A(n11264), .B(n11263), .ZN(
        P2_U3232) );
  INV_X1 U13739 ( .A(n11266), .ZN(n11269) );
  INV_X1 U13740 ( .A(n11267), .ZN(n11268) );
  OAI21_X1 U13741 ( .B1(n11269), .B2(n11268), .A(n11278), .ZN(n12995) );
  XNOR2_X1 U13742 ( .A(n11272), .B(n12995), .ZN(n11270) );
  NAND2_X1 U13743 ( .A1(P3_REG2_REG_15__SCAN_IN), .A2(n11270), .ZN(n12996) );
  OAI21_X1 U13744 ( .B1(P3_REG2_REG_15__SCAN_IN), .B2(n11270), .A(n12996), 
        .ZN(n11286) );
  INV_X1 U13745 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n13741) );
  NOR2_X1 U13746 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13741), .ZN(n12730) );
  AOI21_X1 U13747 ( .B1(n15113), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n12730), 
        .ZN(n11276) );
  NAND2_X1 U13748 ( .A1(n11277), .A2(n11271), .ZN(n13001) );
  OAI21_X1 U13749 ( .B1(n11273), .B2(P3_REG1_REG_15__SCAN_IN), .A(n13002), 
        .ZN(n11274) );
  NAND2_X1 U13750 ( .A1(n13023), .A2(n11274), .ZN(n11275) );
  OAI211_X1 U13751 ( .C1(n15150), .C2(n13010), .A(n11276), .B(n11275), .ZN(
        n11285) );
  MUX2_X1 U13752 ( .A(n11278), .B(n11277), .S(n13037), .Z(n11279) );
  NAND2_X1 U13753 ( .A1(n11280), .A2(n11279), .ZN(n13009) );
  XNOR2_X1 U13754 ( .A(n13009), .B(n13010), .ZN(n11283) );
  INV_X1 U13755 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n11281) );
  INV_X1 U13756 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13328) );
  MUX2_X1 U13757 ( .A(n11281), .B(n13328), .S(n13037), .Z(n11282) );
  NOR2_X1 U13758 ( .A1(n11283), .A2(n11282), .ZN(n13008) );
  AOI211_X1 U13759 ( .C1(n11283), .C2(n11282), .A(n13078), .B(n13008), .ZN(
        n11284) );
  AOI211_X1 U13760 ( .C1(n15154), .C2(n11286), .A(n11285), .B(n11284), .ZN(
        n11287) );
  INV_X1 U13761 ( .A(n11287), .ZN(P3_U3197) );
  MUX2_X1 U13762 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n11907), .Z(n11289) );
  XNOR2_X1 U13763 ( .A(n11289), .B(SI_25_), .ZN(n11330) );
  MUX2_X1 U13764 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n11907), .Z(n11290) );
  NAND2_X1 U13765 ( .A1(n11290), .A2(SI_26_), .ZN(n11291) );
  OAI21_X1 U13766 ( .B1(SI_26_), .B2(n11290), .A(n11291), .ZN(n11424) );
  INV_X1 U13767 ( .A(n11325), .ZN(n11292) );
  NAND2_X1 U13768 ( .A1(n11325), .A2(SI_27_), .ZN(n11293) );
  INV_X1 U13769 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14081) );
  INV_X1 U13770 ( .A(SI_28_), .ZN(n13402) );
  NAND2_X1 U13771 ( .A1(n11295), .A2(n13402), .ZN(n11298) );
  INV_X1 U13772 ( .A(n11295), .ZN(n11296) );
  NAND2_X1 U13773 ( .A1(n11296), .A2(SI_28_), .ZN(n11297) );
  NAND2_X1 U13774 ( .A1(n11298), .A2(n11297), .ZN(n11316) );
  INV_X1 U13775 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n11475) );
  INV_X1 U13776 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14075) );
  MUX2_X1 U13777 ( .A(n11475), .B(n14075), .S(n11907), .Z(n11904) );
  XNOR2_X1 U13778 ( .A(n11904), .B(SI_29_), .ZN(n11902) );
  XNOR2_X1 U13779 ( .A(n11903), .B(n11902), .ZN(n11603) );
  NAND2_X1 U13780 ( .A1(n11603), .A2(n11913), .ZN(n11300) );
  NAND2_X1 U13781 ( .A1(n12116), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n11299) );
  AOI22_X1 U13782 ( .A1(n11459), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n11381), 
        .B2(P1_REG0_REG_29__SCAN_IN), .ZN(n11308) );
  INV_X1 U13783 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n11370) );
  INV_X1 U13784 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14198) );
  NAND2_X1 U13785 ( .A1(n11395), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11394) );
  INV_X1 U13786 ( .A(n11344), .ZN(n11302) );
  NAND2_X1 U13787 ( .A1(n11302), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n11432) );
  INV_X1 U13788 ( .A(n11432), .ZN(n11303) );
  INV_X1 U13789 ( .A(n11434), .ZN(n11305) );
  AND2_X1 U13790 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n11304) );
  NAND2_X1 U13791 ( .A1(n11305), .A2(n11304), .ZN(n11465) );
  INV_X1 U13792 ( .A(n11465), .ZN(n11306) );
  AOI22_X1 U13793 ( .A1(n11320), .A2(P1_REG1_REG_29__SCAN_IN), .B1(n11301), 
        .B2(n11306), .ZN(n11307) );
  NAND2_X1 U13794 ( .A1(n11308), .A2(n11307), .ZN(n14242) );
  XNOR2_X1 U13795 ( .A(n12103), .B(n14242), .ZN(n12157) );
  NAND2_X1 U13796 ( .A1(n11459), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n11315) );
  INV_X1 U13797 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n11309) );
  OR2_X1 U13798 ( .A1(n11921), .A2(n11309), .ZN(n11314) );
  INV_X1 U13799 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n14102) );
  INV_X1 U13800 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n11886) );
  OAI21_X1 U13801 ( .B1(n11434), .B2(n14102), .A(n11886), .ZN(n11310) );
  NAND2_X1 U13802 ( .A1(n11310), .A2(n11465), .ZN(n11890) );
  OR2_X1 U13803 ( .A1(n6575), .A2(n11890), .ZN(n11313) );
  INV_X1 U13804 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n11311) );
  OR2_X1 U13805 ( .A1(n11919), .A2(n11311), .ZN(n11312) );
  NAND4_X1 U13806 ( .A1(n11315), .A2(n11314), .A3(n11313), .A4(n11312), .ZN(
        n14345) );
  NAND2_X1 U13807 ( .A1(n11488), .A2(n11913), .ZN(n11319) );
  NAND2_X1 U13808 ( .A1(n12116), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n11318) );
  NAND2_X1 U13809 ( .A1(n11320), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n11324) );
  INV_X1 U13810 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n13613) );
  OR2_X1 U13811 ( .A1(n11921), .A2(n13613), .ZN(n11323) );
  XNOR2_X1 U13812 ( .A(n11434), .B(n14102), .ZN(n14350) );
  OR2_X1 U13813 ( .A1(n6575), .A2(n14350), .ZN(n11322) );
  INV_X1 U13814 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14351) );
  OR2_X1 U13815 ( .A1(n9229), .A2(n14351), .ZN(n11321) );
  XNOR2_X1 U13816 ( .A(n11325), .B(SI_27_), .ZN(n11326) );
  NAND2_X1 U13817 ( .A1(n11756), .A2(n11913), .ZN(n11329) );
  NAND2_X1 U13818 ( .A1(n12116), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n11328) );
  INV_X1 U13819 ( .A(n14572), .ZN(n14349) );
  XNOR2_X1 U13820 ( .A(n11331), .B(n11330), .ZN(n14085) );
  NAND2_X1 U13821 ( .A1(n14085), .A2(n11913), .ZN(n11333) );
  NAND2_X1 U13822 ( .A1(n12116), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n11332) );
  NAND2_X1 U13823 ( .A1(n11459), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n11341) );
  INV_X1 U13824 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n11334) );
  OR2_X1 U13825 ( .A1(n11921), .A2(n11334), .ZN(n11340) );
  INV_X1 U13826 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n11335) );
  NAND2_X1 U13827 ( .A1(n11344), .A2(n11335), .ZN(n11336) );
  NAND2_X1 U13828 ( .A1(n11432), .A2(n11336), .ZN(n14376) );
  OR2_X1 U13829 ( .A1(n6575), .A2(n14376), .ZN(n11339) );
  INV_X1 U13830 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n11337) );
  OR2_X1 U13831 ( .A1(n11919), .A2(n11337), .ZN(n11338) );
  NAND4_X1 U13832 ( .A1(n11341), .A2(n11340), .A3(n11339), .A4(n11338), .ZN(
        n14392) );
  NAND2_X1 U13833 ( .A1(n11564), .A2(n11913), .ZN(n11343) );
  NAND2_X1 U13834 ( .A1(n12116), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n11342) );
  NAND2_X1 U13835 ( .A1(n11459), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n11349) );
  INV_X1 U13836 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n14665) );
  OR2_X1 U13837 ( .A1(n11921), .A2(n14665), .ZN(n11348) );
  OAI21_X1 U13838 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n11345), .A(n11344), 
        .ZN(n14401) );
  OR2_X1 U13839 ( .A1(n6575), .A2(n14401), .ZN(n11347) );
  INV_X1 U13840 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n14596) );
  OR2_X1 U13841 ( .A1(n11919), .A2(n14596), .ZN(n11346) );
  NAND4_X1 U13842 ( .A1(n11349), .A2(n11348), .A3(n11347), .A4(n11346), .ZN(
        n14244) );
  AND2_X1 U13843 ( .A1(n14647), .A2(n14518), .ZN(n11350) );
  OR2_X1 U13844 ( .A1(n14647), .A2(n14518), .ZN(n11352) );
  NAND2_X1 U13845 ( .A1(n11353), .A2(n11913), .ZN(n11355) );
  AOI22_X1 U13846 ( .A1(n12116), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11366), 
        .B2(n14295), .ZN(n11354) );
  NAND2_X2 U13847 ( .A1(n11355), .A2(n11354), .ZN(n14636) );
  AND2_X1 U13848 ( .A1(n14636), .A2(n14250), .ZN(n11356) );
  NAND2_X1 U13849 ( .A1(n11357), .A2(n11913), .ZN(n11359) );
  AOI22_X1 U13850 ( .A1(n12116), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11366), 
        .B2(n14314), .ZN(n11358) );
  NAND2_X2 U13851 ( .A1(n11359), .A2(n11358), .ZN(n14632) );
  OR2_X1 U13852 ( .A1(n11360), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11361) );
  NAND2_X1 U13853 ( .A1(n11371), .A2(n11361), .ZN(n14503) );
  AOI22_X1 U13854 ( .A1(n11459), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n11381), 
        .B2(P1_REG0_REG_18__SCAN_IN), .ZN(n11364) );
  OR2_X1 U13855 ( .A1(n11919), .A2(n11362), .ZN(n11363) );
  OAI211_X1 U13856 ( .C1(n14503), .C2(n6575), .A(n11364), .B(n11363), .ZN(
        n14249) );
  NOR2_X1 U13857 ( .A1(n14632), .A2(n14249), .ZN(n12042) );
  NAND2_X1 U13858 ( .A1(n14632), .A2(n14249), .ZN(n12041) );
  NAND2_X1 U13859 ( .A1(n11365), .A2(n12041), .ZN(n14477) );
  NAND2_X1 U13860 ( .A1(n11503), .A2(n11913), .ZN(n11369) );
  AOI22_X1 U13861 ( .A1(n12116), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n11367), 
        .B2(n11366), .ZN(n11368) );
  NAND2_X2 U13862 ( .A1(n11369), .A2(n11368), .ZN(n14489) );
  NAND2_X1 U13863 ( .A1(n11371), .A2(n11370), .ZN(n11372) );
  AND2_X1 U13864 ( .A1(n11380), .A2(n11372), .ZN(n14481) );
  NAND2_X1 U13865 ( .A1(n14481), .A2(n11301), .ZN(n11377) );
  INV_X1 U13866 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14311) );
  NAND2_X1 U13867 ( .A1(n8996), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11374) );
  INV_X1 U13868 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14484) );
  OR2_X1 U13869 ( .A1(n9229), .A2(n14484), .ZN(n11373) );
  OAI211_X1 U13870 ( .C1(n14311), .C2(n11919), .A(n11374), .B(n11373), .ZN(
        n11375) );
  INV_X1 U13871 ( .A(n11375), .ZN(n11376) );
  NAND2_X1 U13872 ( .A1(n11377), .A2(n11376), .ZN(n14248) );
  XNOR2_X1 U13873 ( .A(n14489), .B(n14248), .ZN(n12044) );
  NAND2_X1 U13874 ( .A1(n11511), .A2(n11913), .ZN(n11379) );
  NAND2_X1 U13875 ( .A1(n12116), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n11378) );
  AOI21_X1 U13876 ( .B1(n11380), .B2(n14198), .A(n11395), .ZN(n14466) );
  NAND2_X1 U13877 ( .A1(n14466), .A2(n11301), .ZN(n11387) );
  INV_X1 U13878 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n11384) );
  NAND2_X1 U13879 ( .A1(n11459), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n11383) );
  NAND2_X1 U13880 ( .A1(n11381), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11382) );
  OAI211_X1 U13881 ( .C1(n11384), .C2(n11919), .A(n11383), .B(n11382), .ZN(
        n11385) );
  INV_X1 U13882 ( .A(n11385), .ZN(n11386) );
  NAND2_X1 U13883 ( .A1(n11387), .A2(n11386), .ZN(n14247) );
  INV_X1 U13884 ( .A(n14247), .ZN(n11388) );
  NAND2_X1 U13885 ( .A1(n14470), .A2(n11388), .ZN(n11389) );
  NAND2_X1 U13886 ( .A1(n14470), .A2(n14247), .ZN(n11390) );
  NAND2_X1 U13887 ( .A1(n11525), .A2(n11913), .ZN(n11393) );
  OR2_X1 U13888 ( .A1(n11391), .A2(n13655), .ZN(n11392) );
  NAND2_X1 U13889 ( .A1(n8996), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n11400) );
  INV_X1 U13890 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14449) );
  OR2_X1 U13891 ( .A1(n9229), .A2(n14449), .ZN(n11399) );
  OAI21_X1 U13892 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n11395), .A(n11394), 
        .ZN(n14448) );
  OR2_X1 U13893 ( .A1(n6575), .A2(n14448), .ZN(n11398) );
  INV_X1 U13894 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n11396) );
  OR2_X1 U13895 ( .A1(n11919), .A2(n11396), .ZN(n11397) );
  NAND4_X1 U13896 ( .A1(n11400), .A2(n11399), .A3(n11398), .A4(n11397), .ZN(
        n14246) );
  INV_X1 U13897 ( .A(n14246), .ZN(n11448) );
  XNOR2_X1 U13898 ( .A(n14451), .B(n11448), .ZN(n14439) );
  INV_X1 U13899 ( .A(n14439), .ZN(n14444) );
  OR2_X1 U13900 ( .A1(n14451), .A2(n14246), .ZN(n11401) );
  OR2_X1 U13901 ( .A1(n11402), .A2(n11907), .ZN(n11403) );
  NAND2_X1 U13902 ( .A1(n11459), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n11412) );
  INV_X1 U13903 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n11405) );
  OR2_X1 U13904 ( .A1(n11921), .A2(n11405), .ZN(n11411) );
  OAI21_X1 U13905 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n11407), .A(n11406), 
        .ZN(n14433) );
  OR2_X1 U13906 ( .A1(n6575), .A2(n14433), .ZN(n11410) );
  INV_X1 U13907 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n11408) );
  OR2_X1 U13908 ( .A1(n11919), .A2(n11408), .ZN(n11409) );
  INV_X1 U13909 ( .A(n14150), .ZN(n14245) );
  XNOR2_X1 U13910 ( .A(n14606), .B(n14245), .ZN(n14430) );
  NAND2_X1 U13911 ( .A1(n11550), .A2(n11913), .ZN(n11414) );
  NAND2_X1 U13912 ( .A1(n12116), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11413) );
  NAND2_X1 U13913 ( .A1(n11459), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n11422) );
  INV_X1 U13914 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n11415) );
  OR2_X1 U13915 ( .A1(n11921), .A2(n11415), .ZN(n11421) );
  OAI21_X1 U13916 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n11417), .A(n11416), 
        .ZN(n14421) );
  OR2_X1 U13917 ( .A1(n6575), .A2(n14421), .ZN(n11420) );
  INV_X1 U13918 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n11418) );
  OR2_X1 U13919 ( .A1(n11919), .A2(n11418), .ZN(n11419) );
  NAND4_X1 U13920 ( .A1(n11422), .A2(n11421), .A3(n11420), .A4(n11419), .ZN(
        n14393) );
  XNOR2_X1 U13921 ( .A(n14420), .B(n14393), .ZN(n14414) );
  INV_X1 U13922 ( .A(n14414), .ZN(n14410) );
  OR2_X1 U13923 ( .A1(n14420), .A2(n14393), .ZN(n11423) );
  NAND2_X1 U13924 ( .A1(n14409), .A2(n11423), .ZN(n14389) );
  XNOR2_X1 U13925 ( .A(n14403), .B(n14244), .ZN(n14386) );
  INV_X1 U13926 ( .A(n14386), .ZN(n14388) );
  NAND2_X1 U13927 ( .A1(n14389), .A2(n14388), .ZN(n14391) );
  NAND2_X1 U13928 ( .A1(n11425), .A2(n11424), .ZN(n11426) );
  NAND2_X1 U13929 ( .A1(n14082), .A2(n11913), .ZN(n11429) );
  NAND2_X1 U13930 ( .A1(n12116), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n11428) );
  NAND2_X1 U13931 ( .A1(n11459), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n11440) );
  INV_X1 U13932 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n11430) );
  OR2_X1 U13933 ( .A1(n11921), .A2(n11430), .ZN(n11439) );
  INV_X1 U13934 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n11431) );
  NAND2_X1 U13935 ( .A1(n11432), .A2(n11431), .ZN(n11433) );
  NAND2_X1 U13936 ( .A1(n11434), .A2(n11433), .ZN(n14363) );
  OR2_X1 U13937 ( .A1(n6575), .A2(n14363), .ZN(n11438) );
  INV_X1 U13938 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n11436) );
  OR2_X1 U13939 ( .A1(n11919), .A2(n11436), .ZN(n11437) );
  NAND4_X1 U13940 ( .A1(n11440), .A2(n11439), .A3(n11438), .A4(n11437), .ZN(
        n14346) );
  NAND2_X1 U13941 ( .A1(n11862), .A2(n14346), .ZN(n11441) );
  NAND2_X1 U13942 ( .A1(n14578), .A2(n14103), .ZN(n11453) );
  NAND2_X1 U13943 ( .A1(n14566), .A2(n12097), .ZN(n11455) );
  OR2_X1 U13944 ( .A1(n14566), .A2(n12097), .ZN(n11442) );
  NAND2_X1 U13945 ( .A1(n11765), .A2(n12155), .ZN(n11764) );
  OR2_X1 U13946 ( .A1(n14647), .A2(n14251), .ZN(n11443) );
  XNOR2_X1 U13947 ( .A(n14636), .B(n14250), .ZN(n14514) );
  INV_X1 U13948 ( .A(n14250), .ZN(n14493) );
  OR2_X1 U13949 ( .A1(n14636), .A2(n14493), .ZN(n12039) );
  INV_X1 U13950 ( .A(n12042), .ZN(n11445) );
  INV_X1 U13951 ( .A(n14249), .ZN(n14638) );
  INV_X1 U13952 ( .A(n14479), .ZN(n11446) );
  INV_X1 U13953 ( .A(n14248), .ZN(n14494) );
  NAND2_X1 U13954 ( .A1(n14457), .A2(n14461), .ZN(n14456) );
  INV_X1 U13955 ( .A(n14430), .ZN(n11449) );
  INV_X1 U13956 ( .A(n14606), .ZN(n11450) );
  INV_X1 U13957 ( .A(n14393), .ZN(n14188) );
  NAND2_X1 U13958 ( .A1(n14420), .A2(n14188), .ZN(n11451) );
  INV_X1 U13959 ( .A(n14586), .ZN(n11452) );
  INV_X1 U13960 ( .A(n12155), .ZN(n11454) );
  NAND2_X1 U13961 ( .A1(n11758), .A2(n11455), .ZN(n11456) );
  INV_X1 U13962 ( .A(n12103), .ZN(n14559) );
  INV_X1 U13963 ( .A(n14451), .ZN(n14614) );
  NAND2_X1 U13964 ( .A1(n14606), .A2(n14447), .ZN(n14432) );
  NAND2_X1 U13965 ( .A1(n11862), .A2(n11457), .ZN(n14361) );
  AOI21_X1 U13966 ( .B1(n12103), .B2(n11770), .A(n14924), .ZN(n11458) );
  AND2_X2 U13967 ( .A1(n11458), .A2(n14330), .ZN(n14556) );
  NAND2_X1 U13968 ( .A1(n14556), .A2(n14739), .ZN(n11470) );
  INV_X1 U13969 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n11462) );
  NAND2_X1 U13970 ( .A1(n11459), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n11461) );
  NAND2_X1 U13971 ( .A1(n8996), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n11460) );
  OAI211_X1 U13972 ( .C1(n11919), .C2(n11462), .A(n11461), .B(n11460), .ZN(
        n14241) );
  NOR2_X1 U13973 ( .A1(n6663), .A2(n11463), .ZN(n11464) );
  NOR2_X1 U13974 ( .A1(n14637), .A2(n11464), .ZN(n14333) );
  NAND2_X1 U13975 ( .A1(n14241), .A2(n14333), .ZN(n14557) );
  OAI22_X1 U13976 ( .A1(n11466), .A2(n14557), .B1(n11465), .B2(n14541), .ZN(
        n11468) );
  NAND2_X1 U13977 ( .A1(n14345), .A2(n14394), .ZN(n14558) );
  NOR2_X1 U13978 ( .A1(n14743), .A2(n14558), .ZN(n11467) );
  AOI211_X1 U13979 ( .C1(n14743), .C2(P1_REG2_REG_29__SCAN_IN), .A(n11468), 
        .B(n11467), .ZN(n11469) );
  OAI211_X1 U13980 ( .C1(n14559), .C2(n14506), .A(n11470), .B(n11469), .ZN(
        n11471) );
  AOI21_X1 U13981 ( .B1(n14564), .B2(n14480), .A(n11471), .ZN(n11472) );
  OAI21_X1 U13982 ( .B1(n14565), .B2(n14546), .A(n11472), .ZN(P1_U3356) );
  OAI222_X1 U13983 ( .A1(n14088), .A2(n11474), .B1(n14086), .B2(n11512), .C1(
        P2_U3088), .C2(n6629), .ZN(P2_U3307) );
  INV_X1 U13984 ( .A(n11603), .ZN(n14077) );
  OAI222_X1 U13985 ( .A1(n14694), .A2(n14077), .B1(n8693), .B2(P1_U3086), .C1(
        n11475), .C2(n14684), .ZN(P1_U3326) );
  NAND2_X1 U13986 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n11477) );
  INV_X1 U13987 ( .A(n11569), .ZN(n11479) );
  NAND2_X1 U13988 ( .A1(n11479), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n11580) );
  INV_X1 U13989 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13727) );
  INV_X1 U13990 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n11493) );
  INV_X1 U13991 ( .A(n11592), .ZN(n11480) );
  NAND2_X1 U13992 ( .A1(n11480), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n11594) );
  INV_X1 U13993 ( .A(n11594), .ZN(n11481) );
  NAND2_X1 U13994 ( .A1(n11481), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n11629) );
  INV_X1 U13995 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n13466) );
  NAND2_X1 U13996 ( .A1(n11594), .A2(n13466), .ZN(n11482) );
  NAND2_X1 U13997 ( .A1(n11629), .A2(n11482), .ZN(n13602) );
  INV_X1 U13998 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n13950) );
  NAND2_X1 U13999 ( .A1(n11619), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n11484) );
  NAND2_X1 U14000 ( .A1(n10688), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n11483) );
  OAI211_X1 U14001 ( .C1(n13950), .C2(n11609), .A(n11484), .B(n11483), .ZN(
        n11485) );
  INV_X1 U14002 ( .A(n11485), .ZN(n11486) );
  INV_X1 U14003 ( .A(n13534), .ZN(n11602) );
  NAND2_X1 U14004 ( .A1(n11488), .A2(n12393), .ZN(n11490) );
  OR2_X1 U14005 ( .A1(n12400), .A2(n14081), .ZN(n11489) );
  NAND2_X1 U14006 ( .A1(n14082), .A2(n12393), .ZN(n11492) );
  OR2_X1 U14007 ( .A1(n12400), .A2(n14083), .ZN(n11491) );
  NAND2_X1 U14008 ( .A1(n11582), .A2(n11493), .ZN(n11494) );
  NAND2_X1 U14009 ( .A1(n13778), .A2(n6638), .ZN(n11500) );
  INV_X1 U14010 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n11497) );
  NAND2_X1 U14011 ( .A1(n11618), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n11496) );
  NAND2_X1 U14012 ( .A1(n11619), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n11495) );
  OAI211_X1 U14013 ( .C1(n11497), .C2(n11609), .A(n11496), .B(n11495), .ZN(
        n11498) );
  INV_X1 U14014 ( .A(n11498), .ZN(n11499) );
  INV_X1 U14015 ( .A(n13536), .ZN(n11644) );
  OR2_X1 U14016 ( .A1(n14006), .A2(n13445), .ZN(n11501) );
  NAND2_X1 U14017 ( .A1(n11503), .A2(n12393), .ZN(n11507) );
  AOI22_X1 U14018 ( .A1(n11505), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n11504), 
        .B2(n13603), .ZN(n11506) );
  NAND2_X1 U14019 ( .A1(n13899), .A2(n13543), .ZN(n11636) );
  OR2_X1 U14020 ( .A1(n13899), .A2(n13543), .ZN(n11508) );
  NAND2_X1 U14021 ( .A1(n11636), .A2(n11508), .ZN(n13896) );
  INV_X1 U14022 ( .A(n13543), .ZN(n11509) );
  NAND2_X1 U14023 ( .A1(n13899), .A2(n11509), .ZN(n11510) );
  NAND2_X1 U14024 ( .A1(n13889), .A2(n11510), .ZN(n13873) );
  NAND2_X1 U14025 ( .A1(n11511), .A2(n12393), .ZN(n11514) );
  OR2_X1 U14026 ( .A1(n12400), .A2(n11512), .ZN(n11513) );
  INV_X1 U14027 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n11515) );
  NAND2_X1 U14028 ( .A1(n11516), .A2(n11515), .ZN(n11517) );
  NAND2_X1 U14029 ( .A1(n11542), .A2(n11517), .ZN(n13882) );
  OR2_X1 U14030 ( .A1(n13882), .A2(n11606), .ZN(n11522) );
  INV_X1 U14031 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n13997) );
  NAND2_X1 U14032 ( .A1(n11619), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n11519) );
  NAND2_X1 U14033 ( .A1(n11618), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n11518) );
  OAI211_X1 U14034 ( .C1(n13997), .C2(n11609), .A(n11519), .B(n11518), .ZN(
        n11520) );
  INV_X1 U14035 ( .A(n11520), .ZN(n11521) );
  NAND2_X1 U14036 ( .A1(n11522), .A2(n11521), .ZN(n13542) );
  XNOR2_X1 U14037 ( .A(n13881), .B(n13542), .ZN(n13877) );
  INV_X1 U14038 ( .A(n13542), .ZN(n11523) );
  NAND2_X1 U14039 ( .A1(n13881), .A2(n11523), .ZN(n11524) );
  NAND2_X1 U14040 ( .A1(n11525), .A2(n12393), .ZN(n11527) );
  OR2_X1 U14041 ( .A1(n12400), .A2(n13615), .ZN(n11526) );
  XNOR2_X1 U14042 ( .A(n11542), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n13863) );
  NAND2_X1 U14043 ( .A1(n13863), .A2(n6638), .ZN(n11533) );
  INV_X1 U14044 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13731) );
  NAND2_X1 U14045 ( .A1(n12390), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n11530) );
  NAND2_X1 U14046 ( .A1(n11619), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n11529) );
  OAI211_X1 U14047 ( .C1(n9352), .C2(n13731), .A(n11530), .B(n11529), .ZN(
        n11531) );
  INV_X1 U14048 ( .A(n11531), .ZN(n11532) );
  NAND2_X1 U14049 ( .A1(n11533), .A2(n11532), .ZN(n13541) );
  INV_X1 U14050 ( .A(n13541), .ZN(n11691) );
  OR2_X1 U14051 ( .A1(n14050), .A2(n11691), .ZN(n11536) );
  NAND2_X1 U14052 ( .A1(n14050), .A2(n11691), .ZN(n11534) );
  NAND2_X1 U14053 ( .A1(n11536), .A2(n11534), .ZN(n13855) );
  NAND2_X1 U14054 ( .A1(n11537), .A2(n12393), .ZN(n11540) );
  OR2_X1 U14055 ( .A1(n12400), .A2(n11538), .ZN(n11539) );
  INV_X1 U14056 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13474) );
  INV_X1 U14057 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n11541) );
  OAI21_X1 U14058 ( .B1(n11542), .B2(n13474), .A(n11541), .ZN(n11543) );
  NAND2_X1 U14059 ( .A1(n11543), .A2(n11555), .ZN(n13847) );
  OR2_X1 U14060 ( .A1(n13847), .A2(n11606), .ZN(n11548) );
  INV_X1 U14061 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n13986) );
  NAND2_X1 U14062 ( .A1(n11619), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n11545) );
  NAND2_X1 U14063 ( .A1(n11618), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n11544) );
  OAI211_X1 U14064 ( .C1(n13986), .C2(n11609), .A(n11545), .B(n11544), .ZN(
        n11546) );
  INV_X1 U14065 ( .A(n11546), .ZN(n11547) );
  NAND2_X1 U14066 ( .A1(n11548), .A2(n11547), .ZN(n13540) );
  INV_X1 U14067 ( .A(n13540), .ZN(n11694) );
  NAND2_X1 U14068 ( .A1(n13846), .A2(n11694), .ZN(n11549) );
  NAND2_X1 U14069 ( .A1(n11550), .A2(n12393), .ZN(n11553) );
  OR2_X1 U14070 ( .A1(n12400), .A2(n11551), .ZN(n11552) );
  INV_X1 U14071 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n11554) );
  NAND2_X1 U14072 ( .A1(n11555), .A2(n11554), .ZN(n11556) );
  NAND2_X1 U14073 ( .A1(n11569), .A2(n11556), .ZN(n13824) );
  OR2_X1 U14074 ( .A1(n13824), .A2(n11606), .ZN(n11561) );
  INV_X1 U14075 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n13981) );
  NAND2_X1 U14076 ( .A1(n11618), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n11558) );
  NAND2_X1 U14077 ( .A1(n11619), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n11557) );
  OAI211_X1 U14078 ( .C1(n11609), .C2(n13981), .A(n11558), .B(n11557), .ZN(
        n11559) );
  INV_X1 U14079 ( .A(n11559), .ZN(n11560) );
  NAND2_X1 U14080 ( .A1(n11561), .A2(n11560), .ZN(n13539) );
  INV_X1 U14081 ( .A(n13539), .ZN(n11562) );
  OR2_X1 U14082 ( .A1(n13977), .A2(n11562), .ZN(n11563) );
  NAND2_X1 U14083 ( .A1(n13977), .A2(n11562), .ZN(n13803) );
  NAND2_X1 U14084 ( .A1(n11564), .A2(n12393), .ZN(n11567) );
  OR2_X1 U14085 ( .A1(n12400), .A2(n11565), .ZN(n11566) );
  INV_X1 U14086 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n11568) );
  NAND2_X1 U14087 ( .A1(n11569), .A2(n11568), .ZN(n11570) );
  NAND2_X1 U14088 ( .A1(n11580), .A2(n11570), .ZN(n13811) );
  OR2_X1 U14089 ( .A1(n13811), .A2(n11606), .ZN(n11576) );
  INV_X1 U14090 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n11573) );
  NAND2_X1 U14091 ( .A1(n11619), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n11572) );
  NAND2_X1 U14092 ( .A1(n10688), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n11571) );
  OAI211_X1 U14093 ( .C1(n11573), .C2(n11609), .A(n11572), .B(n11571), .ZN(
        n11574) );
  INV_X1 U14094 ( .A(n11574), .ZN(n11575) );
  NAND2_X1 U14095 ( .A1(n11576), .A2(n11575), .ZN(n13538) );
  XNOR2_X1 U14096 ( .A(n13973), .B(n13538), .ZN(n13801) );
  INV_X1 U14097 ( .A(n13538), .ZN(n11729) );
  NAND2_X1 U14098 ( .A1(n13973), .A2(n11729), .ZN(n11577) );
  NAND2_X1 U14099 ( .A1(n13805), .A2(n11577), .ZN(n13786) );
  NAND2_X1 U14100 ( .A1(n14085), .A2(n12393), .ZN(n11579) );
  OR2_X1 U14101 ( .A1(n12400), .A2(n14087), .ZN(n11578) );
  NAND2_X1 U14102 ( .A1(n11580), .A2(n13727), .ZN(n11581) );
  NAND2_X1 U14103 ( .A1(n11582), .A2(n11581), .ZN(n13795) );
  OR2_X1 U14104 ( .A1(n13795), .A2(n11606), .ZN(n11587) );
  INV_X1 U14105 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13969) );
  NAND2_X1 U14106 ( .A1(n11619), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n11584) );
  NAND2_X1 U14107 ( .A1(n11618), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n11583) );
  OAI211_X1 U14108 ( .C1(n13969), .C2(n11609), .A(n11584), .B(n11583), .ZN(
        n11585) );
  INV_X1 U14109 ( .A(n11585), .ZN(n11586) );
  NAND2_X1 U14110 ( .A1(n11587), .A2(n11586), .ZN(n13537) );
  INV_X1 U14111 ( .A(n13537), .ZN(n13513) );
  OR2_X1 U14112 ( .A1(n13964), .A2(n13513), .ZN(n11588) );
  NAND2_X1 U14113 ( .A1(n13964), .A2(n13513), .ZN(n11589) );
  NAND2_X1 U14114 ( .A1(n11756), .A2(n12393), .ZN(n11591) );
  INV_X1 U14115 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n11757) );
  OR2_X1 U14116 ( .A1(n12400), .A2(n11757), .ZN(n11590) );
  INV_X1 U14117 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13430) );
  NAND2_X1 U14118 ( .A1(n11592), .A2(n13430), .ZN(n11593) );
  NAND2_X1 U14119 ( .A1(n11594), .A2(n11593), .ZN(n13763) );
  INV_X1 U14120 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13762) );
  NAND2_X1 U14121 ( .A1(n12390), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n11596) );
  NAND2_X1 U14122 ( .A1(n11619), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n11595) );
  OAI211_X1 U14123 ( .C1(n9352), .C2(n13762), .A(n11596), .B(n11595), .ZN(
        n11597) );
  INV_X1 U14124 ( .A(n11597), .ZN(n11598) );
  INV_X1 U14125 ( .A(n13535), .ZN(n11600) );
  XNOR2_X1 U14126 ( .A(n13954), .B(n11600), .ZN(n13769) );
  INV_X1 U14127 ( .A(n13769), .ZN(n13758) );
  NAND2_X1 U14128 ( .A1(n13608), .A2(n13534), .ZN(n11645) );
  OR2_X1 U14129 ( .A1(n13608), .A2(n13534), .ZN(n11601) );
  NAND2_X1 U14130 ( .A1(n11645), .A2(n11601), .ZN(n13590) );
  NAND2_X1 U14131 ( .A1(n13591), .A2(n13590), .ZN(n13593) );
  OAI21_X1 U14132 ( .B1(n11602), .B2(n13608), .A(n13593), .ZN(n11614) );
  NAND2_X1 U14133 ( .A1(n11603), .A2(n12393), .ZN(n11605) );
  OR2_X1 U14134 ( .A1(n12400), .A2(n14075), .ZN(n11604) );
  OR2_X1 U14135 ( .A1(n11629), .A2(n11606), .ZN(n11613) );
  INV_X1 U14136 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n11610) );
  NAND2_X1 U14137 ( .A1(n11619), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n11608) );
  NAND2_X1 U14138 ( .A1(n10688), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n11607) );
  OAI211_X1 U14139 ( .C1(n11610), .C2(n11609), .A(n11608), .B(n11607), .ZN(
        n11611) );
  INV_X1 U14140 ( .A(n11611), .ZN(n11612) );
  NAND2_X1 U14141 ( .A1(n11613), .A2(n11612), .ZN(n13533) );
  XNOR2_X1 U14142 ( .A(n13944), .B(n13533), .ZN(n12483) );
  NAND2_X1 U14143 ( .A1(n13534), .A2(n13518), .ZN(n11624) );
  INV_X1 U14144 ( .A(P2_B_REG_SCAN_IN), .ZN(n11615) );
  NOR2_X1 U14145 ( .A1(n8501), .A2(n11615), .ZN(n11616) );
  NOR2_X1 U14146 ( .A1(n11617), .A2(n11616), .ZN(n13582) );
  NAND2_X1 U14147 ( .A1(n12390), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n11622) );
  NAND2_X1 U14148 ( .A1(n11618), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n11621) );
  NAND2_X1 U14149 ( .A1(n11619), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n11620) );
  AND3_X1 U14150 ( .A1(n11622), .A2(n11621), .A3(n11620), .ZN(n12405) );
  INV_X1 U14151 ( .A(n12405), .ZN(n13532) );
  INV_X1 U14152 ( .A(n13973), .ZN(n13815) );
  OR2_X2 U14153 ( .A1(n13977), .A2(n13843), .ZN(n13830) );
  NAND2_X1 U14154 ( .A1(n14032), .A2(n11628), .ZN(n13601) );
  AOI211_X1 U14155 ( .C1(n13944), .C2(n13601), .A(n6649), .B(n13586), .ZN(
        n13943) );
  INV_X1 U14156 ( .A(n13944), .ZN(n11632) );
  INV_X1 U14157 ( .A(n11629), .ZN(n11630) );
  AOI22_X1 U14158 ( .A1(n11630), .A2(n15062), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n15075), .ZN(n11631) );
  OAI21_X1 U14159 ( .B1(n11632), .B2(n15069), .A(n11631), .ZN(n11647) );
  INV_X1 U14160 ( .A(n13791), .ZN(n11643) );
  OR2_X1 U14161 ( .A1(n14006), .A2(n13544), .ZN(n11635) );
  INV_X1 U14162 ( .A(n13877), .ZN(n13872) );
  NAND2_X1 U14163 ( .A1(n13878), .A2(n13872), .ZN(n11638) );
  NAND2_X1 U14164 ( .A1(n13881), .A2(n13542), .ZN(n11637) );
  NAND2_X1 U14165 ( .A1(n11638), .A2(n11637), .ZN(n13854) );
  XNOR2_X1 U14166 ( .A(n13846), .B(n13540), .ZN(n13841) );
  NAND2_X1 U14167 ( .A1(n13846), .A2(n13540), .ZN(n11639) );
  INV_X1 U14168 ( .A(n13827), .ZN(n13820) );
  NAND2_X1 U14169 ( .A1(n7199), .A2(n13802), .ZN(n11641) );
  NAND2_X1 U14170 ( .A1(n13973), .A2(n13538), .ZN(n11640) );
  AND2_X1 U14171 ( .A1(n13964), .A2(n13537), .ZN(n11642) );
  NAND2_X1 U14172 ( .A1(n13960), .A2(n13536), .ZN(n12478) );
  NAND2_X1 U14173 ( .A1(n13780), .A2(n11644), .ZN(n12479) );
  INV_X1 U14174 ( .A(n13590), .ZN(n13596) );
  NAND2_X1 U14175 ( .A1(n13597), .A2(n13596), .ZN(n13599) );
  NAND2_X1 U14176 ( .A1(n13599), .A2(n11645), .ZN(n11646) );
  AND2_X1 U14177 ( .A1(n11757), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n11648) );
  INV_X1 U14178 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14685) );
  NAND2_X1 U14179 ( .A1(n14685), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n11650) );
  AND2_X1 U14180 ( .A1(n14681), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n11651) );
  XNOR2_X1 U14181 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n12501) );
  XNOR2_X1 U14182 ( .A(n12503), .B(n12501), .ZN(n13396) );
  NAND2_X1 U14183 ( .A1(n13396), .A2(n12748), .ZN(n11653) );
  INV_X1 U14184 ( .A(SI_29_), .ZN(n13399) );
  OR2_X1 U14185 ( .A1(n6422), .A2(n13399), .ZN(n11652) );
  NAND2_X1 U14186 ( .A1(n11653), .A2(n11652), .ZN(n11669) );
  INV_X1 U14187 ( .A(n12920), .ZN(n11654) );
  AND2_X1 U14188 ( .A1(n12899), .A2(n13111), .ZN(n12902) );
  XNOR2_X1 U14189 ( .A(n14681), .B(P1_DATAO_REG_28__SCAN_IN), .ZN(n11656) );
  NAND2_X1 U14190 ( .A1(n13400), .A2(n12748), .ZN(n11659) );
  OR2_X1 U14191 ( .A1(n6422), .A2(n13402), .ZN(n11658) );
  NAND2_X1 U14192 ( .A1(n13277), .A2(n12569), .ZN(n12904) );
  XOR2_X1 U14193 ( .A(n12949), .B(n12741), .Z(n11901) );
  NAND2_X1 U14194 ( .A1(n13101), .A2(n13111), .ZN(n11660) );
  NAND2_X1 U14195 ( .A1(n11661), .A2(n11660), .ZN(n13088) );
  INV_X1 U14196 ( .A(n13088), .ZN(n11662) );
  NAND2_X1 U14197 ( .A1(n12907), .A2(n12904), .ZN(n12909) );
  NAND2_X1 U14198 ( .A1(n11662), .A2(n12909), .ZN(n13091) );
  OAI21_X1 U14199 ( .B1(n12569), .B2(n13095), .A(n13091), .ZN(n11663) );
  XNOR2_X1 U14200 ( .A(n11663), .B(n12949), .ZN(n11664) );
  NAND2_X1 U14201 ( .A1(n11664), .A2(n14762), .ZN(n11668) );
  NAND2_X1 U14202 ( .A1(n12965), .A2(n15192), .ZN(n11667) );
  NAND2_X1 U14203 ( .A1(n11665), .A2(P3_B_REG_SCAN_IN), .ZN(n11666) );
  NAND2_X1 U14204 ( .A1(n15195), .A2(n11666), .ZN(n13080) );
  AND2_X1 U14205 ( .A1(n11669), .A2(n13311), .ZN(n11898) );
  MUX2_X1 U14206 ( .A(P3_REG1_REG_29__SCAN_IN), .B(n11670), .S(n15240), .Z(
        P3_U3488) );
  XNOR2_X1 U14207 ( .A(n14050), .B(n6627), .ZN(n11692) );
  INV_X1 U14208 ( .A(n11671), .ZN(n11673) );
  NAND2_X1 U14209 ( .A1(n11673), .A2(n11672), .ZN(n11674) );
  XNOR2_X1 U14210 ( .A(n14006), .B(n6627), .ZN(n11676) );
  AND2_X1 U14211 ( .A1(n13544), .A2(n6649), .ZN(n11677) );
  NAND2_X1 U14212 ( .A1(n11676), .A2(n11677), .ZN(n11681) );
  INV_X1 U14213 ( .A(n11676), .ZN(n13446) );
  INV_X1 U14214 ( .A(n11677), .ZN(n11678) );
  NAND2_X1 U14215 ( .A1(n13446), .A2(n11678), .ZN(n11679) );
  NAND2_X1 U14216 ( .A1(n11681), .A2(n11679), .ZN(n13506) );
  XNOR2_X1 U14217 ( .A(n13899), .B(n6627), .ZN(n11683) );
  NAND2_X1 U14218 ( .A1(n13543), .A2(n13845), .ZN(n11684) );
  XNOR2_X1 U14219 ( .A(n11683), .B(n11684), .ZN(n13454) );
  AND2_X1 U14220 ( .A1(n13454), .A2(n11681), .ZN(n11682) );
  INV_X1 U14221 ( .A(n11683), .ZN(n11685) );
  NAND2_X1 U14222 ( .A1(n11685), .A2(n11684), .ZN(n11686) );
  XNOR2_X1 U14223 ( .A(n13881), .B(n13424), .ZN(n11687) );
  NAND2_X1 U14224 ( .A1(n13542), .A2(n13845), .ZN(n11688) );
  NAND2_X1 U14225 ( .A1(n11687), .A2(n11688), .ZN(n13490) );
  INV_X1 U14226 ( .A(n11687), .ZN(n11690) );
  INV_X1 U14227 ( .A(n11688), .ZN(n11689) );
  NAND2_X1 U14228 ( .A1(n11690), .A2(n11689), .ZN(n13489) );
  NOR2_X1 U14229 ( .A1(n11691), .A2(n9326), .ZN(n13471) );
  XNOR2_X1 U14230 ( .A(n13846), .B(n6627), .ZN(n11716) );
  INV_X1 U14231 ( .A(n11695), .ZN(n11696) );
  AOI22_X1 U14232 ( .A1(n11696), .A2(n13527), .B1(n13436), .B2(n13540), .ZN(
        n11701) );
  AOI22_X1 U14233 ( .A1(n13539), .A2(n13517), .B1(n13518), .B2(n13541), .ZN(
        n13836) );
  INV_X1 U14234 ( .A(n13836), .ZN(n11697) );
  AOI22_X1 U14235 ( .A1(n11697), .A2(n13521), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11698) );
  OAI21_X1 U14236 ( .B1(n13847), .B2(n13495), .A(n11698), .ZN(n11699) );
  AOI21_X1 U14237 ( .B1(n13846), .B2(n13510), .A(n11699), .ZN(n11700) );
  OAI21_X1 U14238 ( .B1(n11719), .B2(n11701), .A(n11700), .ZN(P2_U3207) );
  NAND3_X1 U14239 ( .A1(n11702), .A2(n13436), .A3(n13549), .ZN(n11703) );
  OAI21_X1 U14240 ( .B1(n11704), .B2(n13478), .A(n11703), .ZN(n11713) );
  INV_X1 U14241 ( .A(n11705), .ZN(n11712) );
  OAI22_X1 U14242 ( .A1(n13503), .A2(n11707), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11706), .ZN(n11708) );
  AOI21_X1 U14243 ( .B1(n11709), .B2(n13522), .A(n11708), .ZN(n11710) );
  OAI21_X1 U14244 ( .B1(n6959), .B2(n13525), .A(n11710), .ZN(n11711) );
  AOI21_X1 U14245 ( .B1(n11713), .B2(n11712), .A(n11711), .ZN(n11714) );
  OAI21_X1 U14246 ( .B1(n11715), .B2(n13478), .A(n11714), .ZN(P2_U3187) );
  AND2_X1 U14247 ( .A1(n11717), .A2(n11716), .ZN(n11718) );
  XNOR2_X1 U14248 ( .A(n13977), .B(n6627), .ZN(n11721) );
  AND2_X1 U14249 ( .A1(n13539), .A2(n6649), .ZN(n11720) );
  INV_X1 U14250 ( .A(n11721), .ZN(n11722) );
  XNOR2_X1 U14251 ( .A(n13973), .B(n13424), .ZN(n11730) );
  NAND2_X1 U14252 ( .A1(n13538), .A2(n13845), .ZN(n11724) );
  NOR2_X1 U14253 ( .A1(n11730), .A2(n11724), .ZN(n11733) );
  AOI21_X1 U14254 ( .B1(n11730), .B2(n11724), .A(n11733), .ZN(n13481) );
  XNOR2_X1 U14255 ( .A(n13964), .B(n6627), .ZN(n11725) );
  AND2_X1 U14256 ( .A1(n13537), .A2(n6649), .ZN(n11726) );
  NAND2_X1 U14257 ( .A1(n11725), .A2(n11726), .ZN(n13419) );
  INV_X1 U14258 ( .A(n11725), .ZN(n13514) );
  INV_X1 U14259 ( .A(n11726), .ZN(n11727) );
  NAND2_X1 U14260 ( .A1(n13514), .A2(n11727), .ZN(n11728) );
  NAND2_X1 U14261 ( .A1(n13419), .A2(n11728), .ZN(n11734) );
  AOI21_X1 U14262 ( .B1(n13480), .B2(n11734), .A(n13478), .ZN(n11732) );
  NOR3_X1 U14263 ( .A1(n11730), .A2(n11729), .A3(n13512), .ZN(n11731) );
  NOR2_X1 U14264 ( .A1(n11732), .A2(n11731), .ZN(n11741) );
  INV_X1 U14265 ( .A(n11733), .ZN(n11735) );
  NAND2_X1 U14266 ( .A1(n13536), .A2(n13517), .ZN(n11737) );
  NAND2_X1 U14267 ( .A1(n13538), .A2(n13518), .ZN(n11736) );
  NAND2_X1 U14268 ( .A1(n11737), .A2(n11736), .ZN(n13789) );
  AOI22_X1 U14269 ( .A1(n13789), .A2(n13521), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11738) );
  OAI21_X1 U14270 ( .B1(n13795), .B2(n13495), .A(n11738), .ZN(n11739) );
  AOI21_X1 U14271 ( .B1(n13964), .B2(n13510), .A(n11739), .ZN(n11740) );
  OAI21_X1 U14272 ( .B1(n11741), .B2(n13421), .A(n11740), .ZN(P2_U3197) );
  NAND3_X1 U14273 ( .A1(n11742), .A2(n13436), .A3(n13552), .ZN(n11743) );
  OAI21_X1 U14274 ( .B1(n11744), .B2(n13478), .A(n11743), .ZN(n11753) );
  INV_X1 U14275 ( .A(n11745), .ZN(n11752) );
  AOI22_X1 U14276 ( .A1(n13521), .A2(n11746), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11749) );
  NAND2_X1 U14277 ( .A1(n13522), .A2(n11747), .ZN(n11748) );
  OAI211_X1 U14278 ( .C1(n11750), .C2(n13525), .A(n11749), .B(n11748), .ZN(
        n11751) );
  AOI21_X1 U14279 ( .B1(n11753), .B2(n11752), .A(n11751), .ZN(n11754) );
  OAI21_X1 U14280 ( .B1(n11755), .B2(n13478), .A(n11754), .ZN(P2_U3208) );
  INV_X1 U14281 ( .A(n11756), .ZN(n14686) );
  OAI222_X1 U14282 ( .A1(n8501), .A2(P2_U3088), .B1(n14088), .B2(n14686), .C1(
        n11757), .C2(n14086), .ZN(P2_U3300) );
  NAND3_X1 U14283 ( .A1(n7073), .A2(n12155), .A3(n6464), .ZN(n11759) );
  NAND2_X1 U14284 ( .A1(n14243), .A2(n14394), .ZN(n11761) );
  NAND2_X1 U14285 ( .A1(n14242), .A2(n14921), .ZN(n11760) );
  OAI21_X1 U14286 ( .B1(n11765), .B2(n12155), .A(n11764), .ZN(n14570) );
  NAND2_X1 U14287 ( .A1(n14743), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n11766) );
  OAI21_X1 U14288 ( .B1(n14541), .B2(n11890), .A(n11766), .ZN(n11767) );
  AOI21_X1 U14289 ( .B1(n14566), .B2(n14733), .A(n11767), .ZN(n11773) );
  NAND2_X1 U14290 ( .A1(n14566), .A2(n11768), .ZN(n11769) );
  NAND2_X1 U14291 ( .A1(n14567), .A2(n11771), .ZN(n11772) );
  OAI211_X1 U14292 ( .C1(n14570), .C2(n14546), .A(n11773), .B(n11772), .ZN(
        n11774) );
  INV_X1 U14293 ( .A(n11774), .ZN(n11775) );
  OAI21_X1 U14294 ( .B1(n14569), .B2(n14743), .A(n11775), .ZN(P1_U3265) );
  INV_X1 U14295 ( .A(n11776), .ZN(n11778) );
  OAI222_X1 U14296 ( .A1(n9579), .A2(n6925), .B1(n12508), .B2(n11778), .C1(
        n11777), .C2(P3_U3151), .ZN(P3_U3271) );
  OAI22_X1 U14297 ( .A1(n11779), .A2(n8975), .B1(n11780), .B2(n11879), .ZN(
        n11787) );
  INV_X1 U14298 ( .A(n11787), .ZN(n11790) );
  NAND2_X1 U14299 ( .A1(n14119), .A2(n11870), .ZN(n11782) );
  OR2_X1 U14300 ( .A1(n11780), .A2(n8975), .ZN(n11781) );
  NAND2_X1 U14301 ( .A1(n11782), .A2(n11781), .ZN(n11783) );
  XNOR2_X1 U14302 ( .A(n11783), .B(n11881), .ZN(n11788) );
  INV_X1 U14303 ( .A(n11788), .ZN(n11789) );
  XNOR2_X1 U14304 ( .A(n11788), .B(n11787), .ZN(n14111) );
  NAND2_X1 U14305 ( .A1(n14653), .A2(n11870), .ZN(n11792) );
  OR2_X1 U14306 ( .A1(n14113), .A2(n8975), .ZN(n11791) );
  NAND2_X1 U14307 ( .A1(n11792), .A2(n11791), .ZN(n11794) );
  OAI22_X1 U14308 ( .A1(n14240), .A2(n8975), .B1(n14113), .B2(n11879), .ZN(
        n14231) );
  OAI22_X1 U14309 ( .A1(n14647), .A2(n11880), .B1(n14518), .B2(n8975), .ZN(
        n11796) );
  XNOR2_X1 U14310 ( .A(n11796), .B(n11881), .ZN(n11801) );
  OR2_X1 U14311 ( .A1(n14647), .A2(n8975), .ZN(n11798) );
  NAND2_X1 U14312 ( .A1(n14251), .A2(n11874), .ZN(n11797) );
  NAND2_X1 U14313 ( .A1(n11798), .A2(n11797), .ZN(n11800) );
  XNOR2_X1 U14314 ( .A(n11801), .B(n11800), .ZN(n14168) );
  NAND2_X1 U14315 ( .A1(n14636), .A2(n11870), .ZN(n11804) );
  NAND2_X1 U14316 ( .A1(n14250), .A2(n11825), .ZN(n11803) );
  NAND2_X1 U14317 ( .A1(n11804), .A2(n11803), .ZN(n11805) );
  XNOR2_X1 U14318 ( .A(n11805), .B(n11881), .ZN(n11808) );
  AOI22_X1 U14319 ( .A1(n14636), .A2(n6423), .B1(n11874), .B2(n14250), .ZN(
        n11806) );
  XNOR2_X1 U14320 ( .A(n11808), .B(n11806), .ZN(n14177) );
  INV_X1 U14321 ( .A(n11806), .ZN(n11807) );
  INV_X1 U14322 ( .A(n14632), .ZN(n14507) );
  OAI22_X1 U14323 ( .A1(n14507), .A2(n8975), .B1(n14638), .B2(n11879), .ZN(
        n11813) );
  NAND2_X1 U14324 ( .A1(n14632), .A2(n11870), .ZN(n11811) );
  NAND2_X1 U14325 ( .A1(n14249), .A2(n11825), .ZN(n11810) );
  NAND2_X1 U14326 ( .A1(n11811), .A2(n11810), .ZN(n11812) );
  XNOR2_X1 U14327 ( .A(n11812), .B(n11881), .ZN(n11814) );
  XOR2_X1 U14328 ( .A(n11813), .B(n11814), .Z(n14214) );
  NOR2_X1 U14329 ( .A1(n11814), .A2(n11813), .ZN(n11815) );
  NAND2_X1 U14330 ( .A1(n14489), .A2(n11870), .ZN(n11817) );
  NAND2_X1 U14331 ( .A1(n14248), .A2(n11825), .ZN(n11816) );
  NAND2_X1 U14332 ( .A1(n11817), .A2(n11816), .ZN(n11818) );
  XNOR2_X1 U14333 ( .A(n11818), .B(n11881), .ZN(n11822) );
  AND2_X1 U14334 ( .A1(n14248), .A2(n11874), .ZN(n11819) );
  AOI21_X1 U14335 ( .B1(n14489), .B2(n11825), .A(n11819), .ZN(n11820) );
  XNOR2_X1 U14336 ( .A(n11822), .B(n11820), .ZN(n14141) );
  INV_X1 U14337 ( .A(n11820), .ZN(n11821) );
  NAND2_X1 U14338 ( .A1(n11822), .A2(n11821), .ZN(n11823) );
  AND2_X1 U14339 ( .A1(n14247), .A2(n11874), .ZN(n11824) );
  AOI21_X1 U14340 ( .B1(n14470), .B2(n11825), .A(n11824), .ZN(n11828) );
  AOI22_X1 U14341 ( .A1(n14470), .A2(n11870), .B1(n11825), .B2(n14247), .ZN(
        n11826) );
  XNOR2_X1 U14342 ( .A(n11826), .B(n11881), .ZN(n11827) );
  XOR2_X1 U14343 ( .A(n11828), .B(n11827), .Z(n14195) );
  INV_X1 U14344 ( .A(n11827), .ZN(n11830) );
  INV_X1 U14345 ( .A(n11828), .ZN(n11829) );
  NAND2_X1 U14346 ( .A1(n11830), .A2(n11829), .ZN(n11831) );
  AOI22_X1 U14347 ( .A1(n14451), .A2(n11870), .B1(n6423), .B2(n14246), .ZN(
        n11832) );
  XNOR2_X1 U14348 ( .A(n11832), .B(n11881), .ZN(n11834) );
  AOI22_X1 U14349 ( .A1(n14451), .A2(n6423), .B1(n11874), .B2(n14246), .ZN(
        n11833) );
  XNOR2_X1 U14350 ( .A(n11834), .B(n11833), .ZN(n14149) );
  NAND2_X1 U14351 ( .A1(n11834), .A2(n11833), .ZN(n11835) );
  OAI22_X1 U14352 ( .A1(n14606), .A2(n8975), .B1(n14150), .B2(n11879), .ZN(
        n11838) );
  OAI22_X1 U14353 ( .A1(n14606), .A2(n11880), .B1(n14150), .B2(n8975), .ZN(
        n11836) );
  XNOR2_X1 U14354 ( .A(n11836), .B(n11881), .ZN(n11837) );
  XOR2_X1 U14355 ( .A(n11838), .B(n11837), .Z(n14204) );
  INV_X1 U14356 ( .A(n11837), .ZN(n11840) );
  INV_X1 U14357 ( .A(n11838), .ZN(n11839) );
  NAND2_X1 U14358 ( .A1(n11840), .A2(n11839), .ZN(n11841) );
  NAND2_X1 U14359 ( .A1(n14420), .A2(n11870), .ZN(n11843) );
  NAND2_X1 U14360 ( .A1(n14393), .A2(n11825), .ZN(n11842) );
  NAND2_X1 U14361 ( .A1(n11843), .A2(n11842), .ZN(n11844) );
  XNOR2_X1 U14362 ( .A(n11844), .B(n11881), .ZN(n11845) );
  AOI22_X1 U14363 ( .A1(n14420), .A2(n6423), .B1(n11874), .B2(n14393), .ZN(
        n11846) );
  XNOR2_X1 U14364 ( .A(n11845), .B(n11846), .ZN(n14123) );
  INV_X1 U14365 ( .A(n11845), .ZN(n11847) );
  NAND2_X1 U14366 ( .A1(n14403), .A2(n11870), .ZN(n11849) );
  NAND2_X1 U14367 ( .A1(n14244), .A2(n6423), .ZN(n11848) );
  NAND2_X1 U14368 ( .A1(n11849), .A2(n11848), .ZN(n11850) );
  XNOR2_X1 U14369 ( .A(n11850), .B(n11881), .ZN(n11851) );
  AOI22_X1 U14370 ( .A1(n14403), .A2(n6423), .B1(n11874), .B2(n14244), .ZN(
        n11852) );
  XNOR2_X1 U14371 ( .A(n11851), .B(n11852), .ZN(n14184) );
  INV_X1 U14372 ( .A(n11851), .ZN(n11853) );
  NAND2_X1 U14373 ( .A1(n11853), .A2(n11852), .ZN(n11854) );
  NAND2_X1 U14374 ( .A1(n14586), .A2(n11870), .ZN(n11856) );
  NAND2_X1 U14375 ( .A1(n14392), .A2(n6423), .ZN(n11855) );
  NAND2_X1 U14376 ( .A1(n11856), .A2(n11855), .ZN(n11857) );
  XNOR2_X1 U14377 ( .A(n11857), .B(n11881), .ZN(n11858) );
  AOI22_X1 U14378 ( .A1(n14586), .A2(n11825), .B1(n11874), .B2(n14392), .ZN(
        n11859) );
  XNOR2_X1 U14379 ( .A(n11858), .B(n11859), .ZN(n14158) );
  INV_X1 U14380 ( .A(n11858), .ZN(n11860) );
  NAND2_X1 U14381 ( .A1(n11860), .A2(n11859), .ZN(n11861) );
  OAI22_X1 U14382 ( .A1(n11862), .A2(n8975), .B1(n14103), .B2(n11879), .ZN(
        n11867) );
  NAND2_X1 U14383 ( .A1(n14578), .A2(n11870), .ZN(n11864) );
  NAND2_X1 U14384 ( .A1(n14346), .A2(n6423), .ZN(n11863) );
  NAND2_X1 U14385 ( .A1(n11864), .A2(n11863), .ZN(n11865) );
  XNOR2_X1 U14386 ( .A(n11865), .B(n11881), .ZN(n11866) );
  XOR2_X1 U14387 ( .A(n11867), .B(n11866), .Z(n14222) );
  INV_X1 U14388 ( .A(n11866), .ZN(n11869) );
  INV_X1 U14389 ( .A(n11867), .ZN(n11868) );
  NAND2_X1 U14390 ( .A1(n14572), .A2(n11870), .ZN(n11872) );
  NAND2_X1 U14391 ( .A1(n14243), .A2(n11825), .ZN(n11871) );
  NAND2_X1 U14392 ( .A1(n11872), .A2(n11871), .ZN(n11873) );
  XNOR2_X1 U14393 ( .A(n11873), .B(n11881), .ZN(n11876) );
  AOI22_X1 U14394 ( .A1(n14572), .A2(n11825), .B1(n11874), .B2(n14243), .ZN(
        n11877) );
  INV_X1 U14395 ( .A(n11876), .ZN(n11878) );
  OAI22_X1 U14396 ( .A1(n12096), .A2(n8975), .B1(n12097), .B2(n11879), .ZN(
        n11884) );
  OAI22_X1 U14397 ( .A1(n12096), .A2(n11880), .B1(n12097), .B2(n8975), .ZN(
        n11882) );
  XNOR2_X1 U14398 ( .A(n11882), .B(n11881), .ZN(n11883) );
  XOR2_X1 U14399 ( .A(n11884), .B(n11883), .Z(n11885) );
  OAI22_X1 U14400 ( .A1(n14870), .A2(n11887), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11886), .ZN(n11888) );
  AOI21_X1 U14401 ( .B1(n14217), .B2(n14242), .A(n11888), .ZN(n11889) );
  OAI21_X1 U14402 ( .B1(n14883), .B2(n11890), .A(n11889), .ZN(n11891) );
  AOI21_X1 U14403 ( .B1(n14566), .B2(n14879), .A(n11891), .ZN(n11892) );
  OAI21_X1 U14404 ( .B1(n11893), .B2(n14875), .A(n11892), .ZN(P1_U3220) );
  NAND2_X1 U14405 ( .A1(n11894), .A2(n15204), .ZN(n11900) );
  INV_X1 U14406 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n11896) );
  OR2_X1 U14407 ( .A1(n15169), .A2(n11895), .ZN(n13082) );
  OAI21_X1 U14408 ( .B1(n15204), .B2(n11896), .A(n13082), .ZN(n11897) );
  AOI21_X1 U14409 ( .B1(n11898), .B2(n14770), .A(n11897), .ZN(n11899) );
  OAI211_X1 U14410 ( .C1(n11901), .C2(n13207), .A(n11900), .B(n11899), .ZN(
        P3_U3204) );
  NAND2_X1 U14411 ( .A1(n11903), .A2(n11902), .ZN(n11906) );
  NAND2_X1 U14412 ( .A1(n11904), .A2(n13399), .ZN(n11905) );
  NAND2_X1 U14413 ( .A1(n11906), .A2(n11905), .ZN(n12113) );
  MUX2_X1 U14414 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n11907), .Z(n11908) );
  NAND2_X1 U14415 ( .A1(n11908), .A2(SI_30_), .ZN(n11909) );
  OAI21_X1 U14416 ( .B1(SI_30_), .B2(n11908), .A(n11909), .ZN(n12112) );
  MUX2_X1 U14417 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n11907), .Z(n11910) );
  XNOR2_X1 U14418 ( .A(n11910), .B(SI_31_), .ZN(n11911) );
  NAND2_X1 U14419 ( .A1(n14067), .A2(n11913), .ZN(n11915) );
  NAND2_X1 U14420 ( .A1(n12116), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n11914) );
  INV_X4 U14421 ( .A(n12124), .ZN(n12119) );
  NOR2_X1 U14422 ( .A1(n12159), .A2(n12119), .ZN(n12164) );
  INV_X1 U14423 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n11918) );
  NOR2_X1 U14424 ( .A1(n11919), .A2(n11918), .ZN(n11924) );
  INV_X1 U14425 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n13660) );
  NOR2_X1 U14426 ( .A1(n9229), .A2(n13660), .ZN(n11923) );
  INV_X1 U14427 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n11920) );
  NOR2_X1 U14428 ( .A1(n11921), .A2(n11920), .ZN(n11922) );
  NAND2_X1 U14429 ( .A1(n11925), .A2(n6699), .ZN(n11926) );
  NAND2_X1 U14430 ( .A1(n11927), .A2(n11926), .ZN(n11929) );
  NAND2_X1 U14431 ( .A1(n11929), .A2(n11928), .ZN(n12170) );
  NAND2_X1 U14432 ( .A1(n11931), .A2(n11930), .ZN(n12168) );
  NAND2_X1 U14433 ( .A1(n12170), .A2(n12168), .ZN(n12160) );
  NAND2_X1 U14434 ( .A1(n12159), .A2(n12119), .ZN(n12162) );
  NOR2_X1 U14435 ( .A1(n12162), .A2(n14334), .ZN(n11932) );
  AOI211_X1 U14436 ( .C1(n12164), .C2(n14334), .A(n12160), .B(n11932), .ZN(
        n12173) );
  INV_X2 U14437 ( .A(n11933), .ZN(n12076) );
  INV_X1 U14438 ( .A(n12076), .ZN(n12059) );
  MUX2_X1 U14439 ( .A(n12103), .B(n14242), .S(n12059), .Z(n12109) );
  MUX2_X1 U14440 ( .A(n14345), .B(n14566), .S(n12076), .Z(n12099) );
  INV_X1 U14441 ( .A(n12099), .ZN(n12102) );
  NAND2_X1 U14442 ( .A1(n6688), .A2(n14920), .ZN(n11934) );
  NAND2_X1 U14443 ( .A1(n11942), .A2(n11934), .ZN(n11941) );
  OAI211_X1 U14444 ( .C1(n11936), .C2(n11935), .A(n14267), .B(n12076), .ZN(
        n11938) );
  NAND3_X1 U14445 ( .A1(n12076), .A2(n11936), .A3(n11935), .ZN(n11937) );
  OAI211_X1 U14446 ( .C1(n14267), .C2(n11939), .A(n11938), .B(n11937), .ZN(
        n11940) );
  INV_X1 U14447 ( .A(n11942), .ZN(n11943) );
  AND4_X1 U14448 ( .A1(n11957), .A2(n11954), .A3(n9387), .A4(n11945), .ZN(
        n11946) );
  NAND2_X1 U14449 ( .A1(n11951), .A2(n11946), .ZN(n11963) );
  NAND3_X1 U14450 ( .A1(n11957), .A2(n14933), .A3(n12076), .ZN(n11949) );
  NAND3_X1 U14451 ( .A1(n11954), .A2(n11947), .A3(n12119), .ZN(n11948) );
  NAND2_X1 U14452 ( .A1(n11949), .A2(n11948), .ZN(n11950) );
  NAND2_X1 U14453 ( .A1(n11951), .A2(n11950), .ZN(n11962) );
  INV_X1 U14454 ( .A(n11954), .ZN(n11953) );
  OAI211_X1 U14455 ( .C1(n11953), .C2(n11952), .A(n12124), .B(n11957), .ZN(
        n11955) );
  NAND3_X1 U14456 ( .A1(n11958), .A2(n11957), .A3(n11956), .ZN(n11959) );
  NAND2_X1 U14457 ( .A1(n11960), .A2(n11959), .ZN(n11961) );
  NAND3_X1 U14458 ( .A1(n11963), .A2(n11962), .A3(n11961), .ZN(n11969) );
  MUX2_X1 U14459 ( .A(n14263), .B(n11964), .S(n12119), .Z(n11968) );
  OAI21_X1 U14460 ( .B1(n11969), .B2(n11968), .A(n12134), .ZN(n11971) );
  MUX2_X1 U14461 ( .A(n11966), .B(n11965), .S(n12119), .Z(n11967) );
  AOI21_X1 U14462 ( .B1(n11969), .B2(n11968), .A(n11967), .ZN(n11970) );
  AND2_X1 U14463 ( .A1(n14262), .A2(n12076), .ZN(n11974) );
  OAI21_X1 U14464 ( .B1(n14262), .B2(n12124), .A(n11973), .ZN(n11972) );
  OAI21_X1 U14465 ( .B1(n11974), .B2(n11973), .A(n11972), .ZN(n11975) );
  MUX2_X1 U14466 ( .A(n14944), .B(n14261), .S(n12076), .Z(n11978) );
  MUX2_X1 U14467 ( .A(n14944), .B(n14261), .S(n12119), .Z(n11977) );
  MUX2_X1 U14468 ( .A(n14096), .B(n14260), .S(n12119), .Z(n11982) );
  NAND2_X1 U14469 ( .A1(n11981), .A2(n11982), .ZN(n11980) );
  MUX2_X1 U14470 ( .A(n14260), .B(n14096), .S(n12059), .Z(n11979) );
  INV_X1 U14471 ( .A(n11981), .ZN(n11984) );
  INV_X1 U14472 ( .A(n11982), .ZN(n11983) );
  NAND2_X1 U14473 ( .A1(n11984), .A2(n11983), .ZN(n11985) );
  MUX2_X1 U14474 ( .A(n14956), .B(n14259), .S(n12076), .Z(n11987) );
  MUX2_X1 U14475 ( .A(n14956), .B(n14259), .S(n12059), .Z(n11986) );
  MUX2_X1 U14476 ( .A(n14258), .B(n14962), .S(n12076), .Z(n11991) );
  NAND2_X1 U14477 ( .A1(n11990), .A2(n11991), .ZN(n11989) );
  MUX2_X1 U14478 ( .A(n14258), .B(n14962), .S(n12059), .Z(n11988) );
  NAND2_X1 U14479 ( .A1(n11989), .A2(n11988), .ZN(n11995) );
  INV_X1 U14480 ( .A(n11990), .ZN(n11993) );
  INV_X1 U14481 ( .A(n11991), .ZN(n11992) );
  NAND2_X1 U14482 ( .A1(n11993), .A2(n11992), .ZN(n11994) );
  MUX2_X1 U14483 ( .A(n14806), .B(n14257), .S(n12076), .Z(n11997) );
  MUX2_X1 U14484 ( .A(n14806), .B(n14257), .S(n12059), .Z(n11996) );
  MUX2_X1 U14485 ( .A(n14256), .B(n14828), .S(n12076), .Z(n12001) );
  NAND2_X1 U14486 ( .A1(n12000), .A2(n12001), .ZN(n11999) );
  MUX2_X1 U14487 ( .A(n14256), .B(n14828), .S(n12059), .Z(n11998) );
  NAND2_X1 U14488 ( .A1(n11999), .A2(n11998), .ZN(n12005) );
  INV_X1 U14489 ( .A(n12000), .ZN(n12003) );
  INV_X1 U14490 ( .A(n12001), .ZN(n12002) );
  NAND2_X1 U14491 ( .A1(n12003), .A2(n12002), .ZN(n12004) );
  NAND2_X1 U14492 ( .A1(n12005), .A2(n12004), .ZN(n12008) );
  MUX2_X1 U14493 ( .A(n14255), .B(n14734), .S(n12059), .Z(n12009) );
  NAND2_X1 U14494 ( .A1(n12008), .A2(n12009), .ZN(n12007) );
  MUX2_X1 U14495 ( .A(n14255), .B(n14734), .S(n12076), .Z(n12006) );
  NAND2_X1 U14496 ( .A1(n12007), .A2(n12006), .ZN(n12013) );
  INV_X1 U14497 ( .A(n12008), .ZN(n12011) );
  INV_X1 U14498 ( .A(n12009), .ZN(n12010) );
  NAND2_X1 U14499 ( .A1(n12011), .A2(n12010), .ZN(n12012) );
  MUX2_X1 U14500 ( .A(n14835), .B(n14254), .S(n12059), .Z(n12015) );
  INV_X1 U14501 ( .A(n12015), .ZN(n12014) );
  NAND3_X1 U14502 ( .A1(n6450), .A2(n12014), .A3(n12023), .ZN(n12028) );
  NAND2_X1 U14503 ( .A1(n12023), .A2(n14254), .ZN(n12016) );
  MUX2_X1 U14504 ( .A(n12017), .B(n12016), .S(n12076), .Z(n12018) );
  NAND2_X1 U14505 ( .A1(n12024), .A2(n12020), .ZN(n12021) );
  NAND3_X1 U14506 ( .A1(n12021), .A2(n12076), .A3(n12023), .ZN(n12027) );
  NAND2_X1 U14507 ( .A1(n12023), .A2(n12022), .ZN(n12025) );
  NAND3_X1 U14508 ( .A1(n12025), .A2(n12119), .A3(n12024), .ZN(n12026) );
  MUX2_X1 U14509 ( .A(n14518), .B(n14647), .S(n12076), .Z(n12031) );
  NAND2_X1 U14510 ( .A1(n14636), .A2(n14493), .ZN(n12038) );
  MUX2_X1 U14511 ( .A(n12038), .B(n12039), .S(n12059), .Z(n12029) );
  INV_X1 U14512 ( .A(n12030), .ZN(n12037) );
  NAND2_X1 U14513 ( .A1(n12032), .A2(n12031), .ZN(n12035) );
  MUX2_X1 U14514 ( .A(n14251), .B(n14173), .S(n12059), .Z(n12033) );
  NAND2_X1 U14515 ( .A1(n12035), .A2(n12034), .ZN(n12036) );
  MUX2_X1 U14516 ( .A(n12039), .B(n12038), .S(n12059), .Z(n12040) );
  MUX2_X1 U14517 ( .A(n14638), .B(n14507), .S(n12059), .Z(n12043) );
  NAND2_X1 U14518 ( .A1(n14248), .A2(n12124), .ZN(n12046) );
  NAND2_X1 U14519 ( .A1(n14494), .A2(n12119), .ZN(n12045) );
  MUX2_X1 U14520 ( .A(n12046), .B(n12045), .S(n14489), .Z(n12047) );
  MUX2_X1 U14521 ( .A(n14470), .B(n14247), .S(n12059), .Z(n12049) );
  INV_X1 U14522 ( .A(n12049), .ZN(n12051) );
  MUX2_X1 U14523 ( .A(n14247), .B(n14470), .S(n12059), .Z(n12050) );
  NAND2_X1 U14524 ( .A1(n12052), .A2(n12051), .ZN(n12053) );
  MUX2_X1 U14525 ( .A(n14246), .B(n14451), .S(n12059), .Z(n12056) );
  MUX2_X1 U14526 ( .A(n14246), .B(n14451), .S(n12076), .Z(n12055) );
  INV_X1 U14527 ( .A(n12056), .ZN(n12057) );
  MUX2_X1 U14528 ( .A(n14606), .B(n14150), .S(n12059), .Z(n12058) );
  INV_X1 U14529 ( .A(n12058), .ZN(n12061) );
  MUX2_X1 U14530 ( .A(n14150), .B(n14606), .S(n12059), .Z(n12060) );
  AOI21_X1 U14531 ( .B1(n12062), .B2(n12061), .A(n12060), .ZN(n12064) );
  NOR2_X1 U14532 ( .A1(n12062), .A2(n12061), .ZN(n12063) );
  OR2_X1 U14533 ( .A1(n12064), .A2(n12063), .ZN(n12067) );
  MUX2_X1 U14534 ( .A(n14393), .B(n14420), .S(n12119), .Z(n12066) );
  MUX2_X1 U14535 ( .A(n14420), .B(n14393), .S(n12119), .Z(n12065) );
  MUX2_X1 U14536 ( .A(n14403), .B(n14244), .S(n12119), .Z(n12071) );
  MUX2_X1 U14537 ( .A(n14403), .B(n14244), .S(n12076), .Z(n12068) );
  NAND2_X1 U14538 ( .A1(n12069), .A2(n12068), .ZN(n12075) );
  INV_X1 U14539 ( .A(n12070), .ZN(n12073) );
  NAND2_X1 U14540 ( .A1(n12073), .A2(n12072), .ZN(n12074) );
  MUX2_X1 U14541 ( .A(n14586), .B(n14392), .S(n12076), .Z(n12080) );
  NAND2_X1 U14542 ( .A1(n12079), .A2(n12080), .ZN(n12078) );
  MUX2_X1 U14543 ( .A(n14586), .B(n14392), .S(n12119), .Z(n12077) );
  NAND2_X1 U14544 ( .A1(n12078), .A2(n12077), .ZN(n12084) );
  INV_X1 U14545 ( .A(n12079), .ZN(n12082) );
  INV_X1 U14546 ( .A(n12080), .ZN(n12081) );
  NAND2_X1 U14547 ( .A1(n12082), .A2(n12081), .ZN(n12083) );
  MUX2_X1 U14548 ( .A(n14578), .B(n14346), .S(n12119), .Z(n12086) );
  MUX2_X1 U14549 ( .A(n14346), .B(n14578), .S(n12119), .Z(n12085) );
  INV_X1 U14550 ( .A(n12086), .ZN(n12087) );
  MUX2_X1 U14551 ( .A(n14243), .B(n14572), .S(n12119), .Z(n12091) );
  NAND2_X1 U14552 ( .A1(n12090), .A2(n12091), .ZN(n12089) );
  MUX2_X1 U14553 ( .A(n14572), .B(n14243), .S(n12119), .Z(n12088) );
  NAND2_X1 U14554 ( .A1(n12089), .A2(n12088), .ZN(n12095) );
  INV_X1 U14555 ( .A(n12090), .ZN(n12093) );
  INV_X1 U14556 ( .A(n12091), .ZN(n12092) );
  NAND2_X1 U14557 ( .A1(n12093), .A2(n12092), .ZN(n12094) );
  INV_X1 U14558 ( .A(n12100), .ZN(n12101) );
  MUX2_X1 U14559 ( .A(n14242), .B(n12103), .S(n12119), .Z(n12105) );
  NAND2_X1 U14560 ( .A1(n12104), .A2(n12105), .ZN(n12108) );
  INV_X1 U14561 ( .A(n12105), .ZN(n12106) );
  OAI21_X1 U14562 ( .B1(n14334), .B2(n6699), .A(n14241), .ZN(n12111) );
  INV_X1 U14563 ( .A(n12111), .ZN(n12120) );
  NAND2_X1 U14564 ( .A1(n12113), .A2(n12112), .ZN(n12114) );
  NAND2_X1 U14565 ( .A1(n12116), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12117) );
  MUX2_X1 U14566 ( .A(n12120), .B(n14331), .S(n12119), .Z(n12126) );
  INV_X1 U14567 ( .A(n14334), .ZN(n12122) );
  OAI21_X1 U14568 ( .B1(n12122), .B2(n12124), .A(n12121), .ZN(n12123) );
  AOI22_X1 U14569 ( .A1(n14331), .A2(n12076), .B1(n14241), .B2(n12123), .ZN(
        n12125) );
  NAND4_X1 U14570 ( .A1(n12129), .A2(n12130), .A3(n12128), .A4(n12127), .ZN(
        n12132) );
  NOR2_X1 U14571 ( .A1(n12132), .A2(n12131), .ZN(n12135) );
  NAND4_X1 U14572 ( .A1(n12136), .A2(n12135), .A3(n12134), .A4(n12133), .ZN(
        n12137) );
  NOR2_X1 U14573 ( .A1(n12138), .A2(n12137), .ZN(n12141) );
  NAND4_X1 U14574 ( .A1(n12142), .A2(n12141), .A3(n12140), .A4(n12139), .ZN(
        n12143) );
  NOR2_X1 U14575 ( .A1(n12144), .A2(n12143), .ZN(n12146) );
  NAND4_X1 U14576 ( .A1(n14534), .A2(n12147), .A3(n12146), .A4(n12145), .ZN(
        n12148) );
  NOR2_X1 U14577 ( .A1(n12149), .A2(n12148), .ZN(n12150) );
  NAND4_X1 U14578 ( .A1(n14461), .A2(n12150), .A3(n14495), .A4(n14514), .ZN(
        n12151) );
  NOR4_X1 U14579 ( .A1(n14430), .A2(n14478), .A3(n14439), .A4(n12151), .ZN(
        n12152) );
  NAND4_X1 U14580 ( .A1(n14359), .A2(n12152), .A3(n14414), .A4(n14386), .ZN(
        n12154) );
  NOR4_X1 U14581 ( .A1(n12155), .A2(n14344), .A3(n12154), .A4(n12153), .ZN(
        n12158) );
  XNOR2_X1 U14582 ( .A(n14331), .B(n14241), .ZN(n12156) );
  NOR3_X1 U14583 ( .A1(n14552), .A2(n14334), .A3(n12160), .ZN(n12163) );
  NOR3_X1 U14584 ( .A1(n12162), .A2(n14334), .A3(n12170), .ZN(n12161) );
  AOI21_X1 U14585 ( .B1(n12163), .B2(n12162), .A(n12161), .ZN(n12167) );
  XOR2_X1 U14586 ( .A(n12170), .B(n12164), .Z(n12165) );
  NAND4_X1 U14587 ( .A1(n12165), .A2(n14552), .A3(n14334), .A4(n12168), .ZN(
        n12166) );
  OAI211_X1 U14588 ( .C1(n12169), .C2(n12168), .A(n12167), .B(n12166), .ZN(
        n12172) );
  NAND3_X1 U14589 ( .A1(n12175), .A2(n12174), .A3(n14394), .ZN(n12176) );
  OAI211_X1 U14590 ( .C1(n8784), .C2(n12178), .A(n12176), .B(P1_B_REG_SCAN_IN), 
        .ZN(n12177) );
  INV_X1 U14591 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12504) );
  NAND2_X1 U14592 ( .A1(n12184), .A2(n12186), .ZN(n12182) );
  OAI211_X1 U14593 ( .C1(n12183), .C2(n12432), .A(n12182), .B(n12185), .ZN(
        n12190) );
  OAI21_X1 U14594 ( .B1(n12185), .B2(n12444), .A(n12184), .ZN(n12188) );
  INV_X1 U14595 ( .A(n12186), .ZN(n12187) );
  NAND2_X1 U14596 ( .A1(n12188), .A2(n12187), .ZN(n12189) );
  NAND2_X1 U14597 ( .A1(n12432), .A2(n13926), .ZN(n12192) );
  AND2_X1 U14598 ( .A1(n12192), .A2(n12191), .ZN(n12196) );
  NAND2_X1 U14599 ( .A1(n12432), .A2(n13561), .ZN(n12193) );
  OAI21_X1 U14600 ( .B1(n12194), .B2(n12432), .A(n12193), .ZN(n12195) );
  NAND2_X1 U14601 ( .A1(n12197), .A2(n12196), .ZN(n12198) );
  INV_X2 U14602 ( .A(n12432), .ZN(n12397) );
  NAND2_X1 U14603 ( .A1(n12397), .A2(n13916), .ZN(n12201) );
  NAND2_X1 U14605 ( .A1(n12432), .A2(n13560), .ZN(n12200) );
  NAND2_X1 U14606 ( .A1(n12201), .A2(n12200), .ZN(n12207) );
  NAND2_X1 U14607 ( .A1(n12206), .A2(n12207), .ZN(n12205) );
  NAND2_X1 U14608 ( .A1(n13916), .A2(n12432), .ZN(n12202) );
  NAND2_X1 U14609 ( .A1(n12205), .A2(n12204), .ZN(n12211) );
  INV_X1 U14610 ( .A(n12206), .ZN(n12209) );
  INV_X1 U14611 ( .A(n12207), .ZN(n12208) );
  NAND2_X1 U14612 ( .A1(n12209), .A2(n12208), .ZN(n12210) );
  NAND2_X1 U14613 ( .A1(n12408), .A2(n13559), .ZN(n12213) );
  NAND2_X1 U14614 ( .A1(n13908), .A2(n12412), .ZN(n12212) );
  NAND2_X1 U14615 ( .A1(n12213), .A2(n12212), .ZN(n12216) );
  AOI22_X1 U14616 ( .A1(n12397), .A2(n13908), .B1(n12412), .B2(n13559), .ZN(
        n12215) );
  NAND2_X1 U14617 ( .A1(n15089), .A2(n12397), .ZN(n12219) );
  NAND2_X1 U14618 ( .A1(n12412), .A2(n13558), .ZN(n12218) );
  NAND2_X1 U14619 ( .A1(n12219), .A2(n12218), .ZN(n12221) );
  AOI22_X1 U14620 ( .A1(n15089), .A2(n12412), .B1(n12408), .B2(n13558), .ZN(
        n12220) );
  INV_X2 U14621 ( .A(n12397), .ZN(n12403) );
  NAND2_X1 U14622 ( .A1(n12227), .A2(n12403), .ZN(n12225) );
  NAND2_X1 U14623 ( .A1(n12408), .A2(n13557), .ZN(n12224) );
  NAND2_X1 U14624 ( .A1(n12225), .A2(n12224), .ZN(n12226) );
  AOI22_X1 U14625 ( .A1(n12227), .A2(n12408), .B1(n13557), .B2(n12403), .ZN(
        n12228) );
  NAND2_X1 U14626 ( .A1(n15097), .A2(n12408), .ZN(n12230) );
  NAND2_X1 U14627 ( .A1(n12403), .A2(n13556), .ZN(n12229) );
  NAND2_X1 U14628 ( .A1(n12230), .A2(n12229), .ZN(n12235) );
  NAND2_X1 U14629 ( .A1(n12234), .A2(n12235), .ZN(n12233) );
  NAND2_X1 U14630 ( .A1(n15097), .A2(n12403), .ZN(n12231) );
  OAI21_X1 U14631 ( .B1(n13404), .B2(n12432), .A(n12231), .ZN(n12232) );
  NAND2_X1 U14632 ( .A1(n12233), .A2(n12232), .ZN(n12239) );
  INV_X1 U14633 ( .A(n12234), .ZN(n12237) );
  INV_X1 U14634 ( .A(n12235), .ZN(n12236) );
  NAND2_X1 U14635 ( .A1(n12237), .A2(n12236), .ZN(n12238) );
  NAND2_X1 U14636 ( .A1(n13414), .A2(n12403), .ZN(n12241) );
  NAND2_X1 U14637 ( .A1(n12408), .A2(n13555), .ZN(n12240) );
  AOI22_X1 U14638 ( .A1(n13414), .A2(n12408), .B1(n13555), .B2(n12403), .ZN(
        n12242) );
  NAND2_X1 U14639 ( .A1(n12245), .A2(n12408), .ZN(n12244) );
  NAND2_X1 U14640 ( .A1(n12403), .A2(n13554), .ZN(n12243) );
  NAND2_X1 U14641 ( .A1(n12244), .A2(n12243), .ZN(n12249) );
  NAND2_X1 U14642 ( .A1(n12250), .A2(n12249), .ZN(n12248) );
  AOI22_X1 U14643 ( .A1(n12245), .A2(n12403), .B1(n12408), .B2(n13554), .ZN(
        n12246) );
  NAND2_X1 U14644 ( .A1(n12248), .A2(n12247), .ZN(n12252) );
  INV_X1 U14645 ( .A(n12258), .ZN(n12256) );
  NAND2_X1 U14646 ( .A1(n12259), .A2(n12403), .ZN(n12254) );
  NAND2_X1 U14647 ( .A1(n12408), .A2(n13553), .ZN(n12253) );
  NAND2_X1 U14648 ( .A1(n12254), .A2(n12253), .ZN(n12257) );
  INV_X1 U14649 ( .A(n12257), .ZN(n12255) );
  NAND2_X1 U14650 ( .A1(n12256), .A2(n12255), .ZN(n12265) );
  NAND2_X1 U14651 ( .A1(n12259), .A2(n12408), .ZN(n12260) );
  OAI21_X1 U14652 ( .B1(n12261), .B2(n12408), .A(n12260), .ZN(n12262) );
  NAND2_X1 U14653 ( .A1(n12263), .A2(n12262), .ZN(n12264) );
  NAND2_X1 U14654 ( .A1(n12268), .A2(n12408), .ZN(n12267) );
  NAND2_X1 U14655 ( .A1(n12403), .A2(n13552), .ZN(n12266) );
  AOI22_X1 U14656 ( .A1(n12268), .A2(n12403), .B1(n12408), .B2(n13552), .ZN(
        n12269) );
  NAND2_X1 U14657 ( .A1(n6651), .A2(n12403), .ZN(n12272) );
  NAND2_X1 U14658 ( .A1(n12408), .A2(n13551), .ZN(n12271) );
  NAND2_X1 U14659 ( .A1(n6651), .A2(n12408), .ZN(n12275) );
  NAND2_X1 U14660 ( .A1(n12403), .A2(n13551), .ZN(n12274) );
  NAND2_X1 U14661 ( .A1(n12275), .A2(n12274), .ZN(n12276) );
  NAND2_X1 U14662 ( .A1(n12277), .A2(n12276), .ZN(n12278) );
  NAND2_X1 U14663 ( .A1(n12278), .A2(n7426), .ZN(n12284) );
  NAND2_X1 U14664 ( .A1(n6604), .A2(n12408), .ZN(n12280) );
  NAND2_X1 U14665 ( .A1(n12403), .A2(n13550), .ZN(n12279) );
  NAND2_X1 U14666 ( .A1(n12280), .A2(n12279), .ZN(n12283) );
  AOI22_X1 U14667 ( .A1(n6604), .A2(n12403), .B1(n12408), .B2(n13550), .ZN(
        n12282) );
  NAND2_X1 U14668 ( .A1(n14017), .A2(n12403), .ZN(n12288) );
  NAND2_X1 U14669 ( .A1(n12408), .A2(n13549), .ZN(n12287) );
  NAND2_X1 U14670 ( .A1(n14017), .A2(n12408), .ZN(n12289) );
  OAI21_X1 U14671 ( .B1(n12290), .B2(n12397), .A(n12289), .ZN(n12291) );
  NAND2_X1 U14672 ( .A1(n6593), .A2(n12408), .ZN(n12293) );
  NAND2_X1 U14673 ( .A1(n13548), .A2(n12403), .ZN(n12292) );
  NAND2_X1 U14674 ( .A1(n12293), .A2(n12292), .ZN(n12296) );
  AOI22_X1 U14675 ( .A1(n6593), .A2(n12403), .B1(n12408), .B2(n13548), .ZN(
        n12295) );
  NAND2_X1 U14676 ( .A1(n12300), .A2(n12403), .ZN(n12299) );
  NAND2_X1 U14677 ( .A1(n13547), .A2(n12408), .ZN(n12298) );
  NAND2_X1 U14678 ( .A1(n12299), .A2(n12298), .ZN(n12302) );
  NOR2_X1 U14679 ( .A1(n12303), .A2(n12302), .ZN(n12304) );
  NAND2_X1 U14680 ( .A1(n12308), .A2(n12408), .ZN(n12307) );
  NAND2_X1 U14681 ( .A1(n13546), .A2(n12403), .ZN(n12306) );
  NAND2_X1 U14682 ( .A1(n12308), .A2(n12403), .ZN(n12309) );
  OAI21_X1 U14683 ( .B1(n12310), .B2(n12432), .A(n12309), .ZN(n12311) );
  NAND2_X1 U14684 ( .A1(n12314), .A2(n12403), .ZN(n12313) );
  NAND2_X1 U14685 ( .A1(n13545), .A2(n12408), .ZN(n12312) );
  NAND2_X1 U14686 ( .A1(n12313), .A2(n12312), .ZN(n12317) );
  INV_X1 U14687 ( .A(n12316), .ZN(n12319) );
  NAND2_X1 U14688 ( .A1(n14006), .A2(n12408), .ZN(n12321) );
  NAND2_X1 U14689 ( .A1(n13544), .A2(n12403), .ZN(n12320) );
  NAND2_X1 U14690 ( .A1(n12321), .A2(n12320), .ZN(n12326) );
  NAND2_X1 U14691 ( .A1(n14006), .A2(n12403), .ZN(n12322) );
  NAND2_X1 U14692 ( .A1(n12324), .A2(n12323), .ZN(n12330) );
  INV_X1 U14693 ( .A(n12325), .ZN(n12328) );
  INV_X1 U14694 ( .A(n12326), .ZN(n12327) );
  NAND2_X1 U14695 ( .A1(n12328), .A2(n12327), .ZN(n12329) );
  NAND2_X1 U14696 ( .A1(n13899), .A2(n12403), .ZN(n12332) );
  NAND2_X1 U14697 ( .A1(n13543), .A2(n12408), .ZN(n12331) );
  AOI22_X1 U14698 ( .A1(n13899), .A2(n12408), .B1(n13543), .B2(n12403), .ZN(
        n12333) );
  NAND2_X1 U14699 ( .A1(n13881), .A2(n12408), .ZN(n12335) );
  NAND2_X1 U14700 ( .A1(n13542), .A2(n12403), .ZN(n12334) );
  NAND2_X1 U14701 ( .A1(n12335), .A2(n12334), .ZN(n12338) );
  AOI22_X1 U14702 ( .A1(n13881), .A2(n12403), .B1(n12408), .B2(n13542), .ZN(
        n12336) );
  NAND2_X1 U14703 ( .A1(n14050), .A2(n12403), .ZN(n12341) );
  NAND2_X1 U14704 ( .A1(n13541), .A2(n12408), .ZN(n12340) );
  NAND2_X1 U14705 ( .A1(n14050), .A2(n12408), .ZN(n12343) );
  NAND2_X1 U14706 ( .A1(n13541), .A2(n12412), .ZN(n12342) );
  NAND2_X1 U14707 ( .A1(n12343), .A2(n12342), .ZN(n12344) );
  NAND2_X1 U14708 ( .A1(n13846), .A2(n12408), .ZN(n12346) );
  NAND2_X1 U14709 ( .A1(n13540), .A2(n12403), .ZN(n12345) );
  NAND2_X1 U14710 ( .A1(n12346), .A2(n12345), .ZN(n12348) );
  AOI22_X1 U14711 ( .A1(n13846), .A2(n12412), .B1(n12408), .B2(n13540), .ZN(
        n12347) );
  NAND2_X1 U14712 ( .A1(n13977), .A2(n12403), .ZN(n12352) );
  NAND2_X1 U14713 ( .A1(n13539), .A2(n12408), .ZN(n12351) );
  NAND2_X1 U14714 ( .A1(n12352), .A2(n12351), .ZN(n12353) );
  NAND2_X1 U14715 ( .A1(n12354), .A2(n12353), .ZN(n12358) );
  NAND2_X1 U14716 ( .A1(n13977), .A2(n12397), .ZN(n12356) );
  NAND2_X1 U14717 ( .A1(n13539), .A2(n12412), .ZN(n12355) );
  NAND2_X1 U14718 ( .A1(n12356), .A2(n12355), .ZN(n12357) );
  NAND2_X1 U14719 ( .A1(n13973), .A2(n12397), .ZN(n12360) );
  NAND2_X1 U14720 ( .A1(n13538), .A2(n12412), .ZN(n12359) );
  AOI22_X1 U14721 ( .A1(n13973), .A2(n12412), .B1(n12408), .B2(n13538), .ZN(
        n12361) );
  AND2_X1 U14722 ( .A1(n13536), .A2(n12408), .ZN(n12362) );
  AOI21_X1 U14723 ( .B1(n13960), .B2(n12412), .A(n12362), .ZN(n12375) );
  NAND2_X1 U14724 ( .A1(n13960), .A2(n12408), .ZN(n12364) );
  NAND2_X1 U14725 ( .A1(n13536), .A2(n12412), .ZN(n12363) );
  NAND2_X1 U14726 ( .A1(n12364), .A2(n12363), .ZN(n12374) );
  NAND2_X1 U14727 ( .A1(n12375), .A2(n12374), .ZN(n12379) );
  AND2_X1 U14728 ( .A1(n13537), .A2(n12403), .ZN(n12365) );
  AOI21_X1 U14729 ( .B1(n13964), .B2(n12397), .A(n12365), .ZN(n12373) );
  NAND2_X1 U14730 ( .A1(n13964), .A2(n12403), .ZN(n12367) );
  NAND2_X1 U14731 ( .A1(n13537), .A2(n12408), .ZN(n12366) );
  NAND2_X1 U14732 ( .A1(n12367), .A2(n12366), .ZN(n12372) );
  AND2_X1 U14733 ( .A1(n13535), .A2(n12403), .ZN(n12369) );
  AOI21_X1 U14734 ( .B1(n13954), .B2(n12408), .A(n12369), .ZN(n12386) );
  NAND2_X1 U14735 ( .A1(n13954), .A2(n12403), .ZN(n12371) );
  NAND2_X1 U14736 ( .A1(n13535), .A2(n12397), .ZN(n12370) );
  NAND2_X1 U14737 ( .A1(n12371), .A2(n12370), .ZN(n12385) );
  NAND2_X1 U14738 ( .A1(n12386), .A2(n12385), .ZN(n12381) );
  AND2_X1 U14739 ( .A1(n12373), .A2(n12372), .ZN(n12378) );
  INV_X1 U14740 ( .A(n12374), .ZN(n12377) );
  INV_X1 U14741 ( .A(n12375), .ZN(n12376) );
  AOI22_X1 U14742 ( .A1(n12379), .A2(n12378), .B1(n12377), .B2(n12376), .ZN(
        n12380) );
  AND2_X1 U14743 ( .A1(n13534), .A2(n12408), .ZN(n12382) );
  AOI21_X1 U14744 ( .B1(n13608), .B2(n12403), .A(n12382), .ZN(n12421) );
  NAND2_X1 U14745 ( .A1(n13608), .A2(n12397), .ZN(n12384) );
  NAND2_X1 U14746 ( .A1(n13534), .A2(n12412), .ZN(n12383) );
  NAND2_X1 U14747 ( .A1(n12384), .A2(n12383), .ZN(n12420) );
  INV_X1 U14748 ( .A(n12385), .ZN(n12388) );
  INV_X1 U14749 ( .A(n12386), .ZN(n12387) );
  AOI22_X1 U14750 ( .A1(n12421), .A2(n12420), .B1(n12388), .B2(n12387), .ZN(
        n12389) );
  INV_X1 U14751 ( .A(n12389), .ZN(n12418) );
  INV_X1 U14752 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n14022) );
  NAND2_X1 U14753 ( .A1(n12390), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n12392) );
  NAND2_X1 U14754 ( .A1(n10688), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n12391) );
  OAI211_X1 U14755 ( .C1(n8942), .C2(n14022), .A(n12392), .B(n12391), .ZN(
        n13581) );
  NAND2_X1 U14756 ( .A1(n14067), .A2(n12393), .ZN(n12396) );
  INV_X1 U14757 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12394) );
  OR2_X1 U14758 ( .A1(n12400), .A2(n12394), .ZN(n12395) );
  MUX2_X1 U14759 ( .A(n13581), .B(n12397), .S(n13579), .Z(n12398) );
  NAND2_X1 U14760 ( .A1(n12408), .A2(n13581), .ZN(n12431) );
  NAND2_X1 U14761 ( .A1(n12398), .A2(n12431), .ZN(n12416) );
  INV_X1 U14762 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n14072) );
  OR2_X1 U14763 ( .A1(n12400), .A2(n14072), .ZN(n12401) );
  NAND2_X1 U14764 ( .A1(n12403), .A2(n13581), .ZN(n12433) );
  NAND2_X1 U14765 ( .A1(n12489), .A2(n12498), .ZN(n12440) );
  AND2_X1 U14766 ( .A1(n12404), .A2(n12440), .ZN(n12406) );
  AOI21_X1 U14767 ( .B1(n12433), .B2(n12406), .A(n12405), .ZN(n12407) );
  AOI21_X1 U14768 ( .B1(n13940), .B2(n12397), .A(n12407), .ZN(n12428) );
  NAND2_X1 U14769 ( .A1(n13940), .A2(n12412), .ZN(n12410) );
  NAND2_X1 U14770 ( .A1(n12408), .A2(n13532), .ZN(n12409) );
  NAND2_X1 U14771 ( .A1(n12410), .A2(n12409), .ZN(n12427) );
  AND2_X1 U14772 ( .A1(n13533), .A2(n12412), .ZN(n12411) );
  AOI21_X1 U14773 ( .B1(n13944), .B2(n12397), .A(n12411), .ZN(n12425) );
  NAND2_X1 U14774 ( .A1(n13944), .A2(n12412), .ZN(n12414) );
  NAND2_X1 U14775 ( .A1(n13533), .A2(n12397), .ZN(n12413) );
  NAND2_X1 U14776 ( .A1(n12414), .A2(n12413), .ZN(n12424) );
  OAI22_X1 U14777 ( .A1(n12428), .A2(n12427), .B1(n12425), .B2(n12424), .ZN(
        n12415) );
  NAND2_X1 U14778 ( .A1(n12416), .A2(n12415), .ZN(n12430) );
  XNOR2_X1 U14779 ( .A(n13579), .B(n13581), .ZN(n12484) );
  INV_X1 U14780 ( .A(n12420), .ZN(n12423) );
  INV_X1 U14781 ( .A(n12421), .ZN(n12422) );
  AOI22_X1 U14782 ( .A1(n12425), .A2(n12424), .B1(n12423), .B2(n12422), .ZN(
        n12426) );
  NAND2_X1 U14783 ( .A1(n12484), .A2(n12426), .ZN(n12429) );
  AOI22_X1 U14784 ( .A1(n12430), .A2(n12429), .B1(n12428), .B2(n12427), .ZN(
        n12437) );
  INV_X1 U14785 ( .A(n12431), .ZN(n12435) );
  AND2_X1 U14786 ( .A1(n12433), .A2(n12432), .ZN(n12434) );
  MUX2_X1 U14787 ( .A(n12435), .B(n12434), .S(n13579), .Z(n12436) );
  NAND3_X1 U14788 ( .A1(n12449), .A2(n12488), .A3(n13603), .ZN(n12439) );
  NAND2_X1 U14789 ( .A1(n12441), .A2(n13574), .ZN(n12442) );
  OAI211_X1 U14790 ( .C1(n12444), .C2(n12498), .A(n12443), .B(n12442), .ZN(
        n12445) );
  NAND2_X1 U14791 ( .A1(n12490), .A2(n12445), .ZN(n12446) );
  OAI21_X1 U14792 ( .B1(n12490), .B2(n6560), .A(n12446), .ZN(n12493) );
  XOR2_X1 U14793 ( .A(n13532), .B(n13940), .Z(n12482) );
  NAND4_X1 U14794 ( .A1(n12450), .A2(n12449), .A3(n12448), .A4(n12447), .ZN(
        n12452) );
  NOR2_X1 U14795 ( .A1(n12452), .A2(n12451), .ZN(n12455) );
  NAND4_X1 U14796 ( .A1(n12456), .A2(n12455), .A3(n12454), .A4(n12453), .ZN(
        n12457) );
  NOR2_X1 U14797 ( .A1(n12458), .A2(n12457), .ZN(n12461) );
  NAND4_X1 U14798 ( .A1(n12462), .A2(n12461), .A3(n12460), .A4(n12459), .ZN(
        n12463) );
  NOR2_X1 U14799 ( .A1(n12464), .A2(n12463), .ZN(n12467) );
  NAND4_X1 U14800 ( .A1(n12468), .A2(n12467), .A3(n12466), .A4(n12465), .ZN(
        n12469) );
  OR3_X1 U14801 ( .A1(n12471), .A2(n12470), .A3(n12469), .ZN(n12472) );
  NOR2_X1 U14802 ( .A1(n12473), .A2(n12472), .ZN(n12474) );
  NAND3_X1 U14803 ( .A1(n13877), .A2(n13896), .A3(n12474), .ZN(n12476) );
  NOR3_X1 U14804 ( .A1(n13855), .A2(n12476), .A3(n12475), .ZN(n12477) );
  AND4_X1 U14805 ( .A1(n13801), .A2(n13827), .A3(n12477), .A4(n13841), .ZN(
        n12480) );
  NAND2_X1 U14806 ( .A1(n12479), .A2(n12478), .ZN(n13781) );
  NAND4_X1 U14807 ( .A1(n13590), .A2(n13791), .A3(n12480), .A4(n13781), .ZN(
        n12481) );
  NOR3_X1 U14808 ( .A1(n12482), .A2(n13769), .A3(n12481), .ZN(n12485) );
  NAND3_X1 U14809 ( .A1(n12485), .A2(n12484), .A3(n12483), .ZN(n12486) );
  XOR2_X1 U14810 ( .A(n13603), .B(n12486), .Z(n12487) );
  OAI21_X1 U14811 ( .B1(n12493), .B2(n12492), .A(n12491), .ZN(n12500) );
  INV_X1 U14812 ( .A(n8501), .ZN(n12495) );
  NAND4_X1 U14813 ( .A1(n15087), .A2(n12495), .A3(n12494), .A4(n13518), .ZN(
        n12496) );
  OAI211_X1 U14814 ( .C1(n12498), .C2(n12497), .A(n12496), .B(P2_B_REG_SCAN_IN), .ZN(n12499) );
  NAND2_X1 U14815 ( .A1(n12500), .A2(n12499), .ZN(P2_U3328) );
  INV_X1 U14816 ( .A(SI_30_), .ZN(n12750) );
  INV_X1 U14817 ( .A(n12501), .ZN(n12502) );
  OAI22_X1 U14818 ( .A1(n12503), .A2(n12502), .B1(P2_DATAO_REG_29__SCAN_IN), 
        .B2(n14075), .ZN(n12743) );
  NAND2_X1 U14819 ( .A1(n14072), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12744) );
  NAND2_X1 U14820 ( .A1(n12504), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12505) );
  NAND2_X1 U14821 ( .A1(n12744), .A2(n12505), .ZN(n12742) );
  XNOR2_X1 U14822 ( .A(n12743), .B(n12742), .ZN(n12749) );
  INV_X1 U14823 ( .A(n12749), .ZN(n12507) );
  OAI222_X1 U14824 ( .A1(n9579), .A2(n12750), .B1(n12508), .B2(n12507), .C1(
        n12506), .C2(P3_U3151), .ZN(P3_U3265) );
  INV_X1 U14825 ( .A(n12509), .ZN(n12510) );
  OAI222_X1 U14826 ( .A1(n9579), .A2(n12511), .B1(n12508), .B2(n12510), .C1(
        n13037), .C2(P3_U3151), .ZN(P3_U3268) );
  OR2_X1 U14827 ( .A1(n12512), .A2(n12970), .ZN(n12513) );
  XNOR2_X1 U14828 ( .A(n12614), .B(n15227), .ZN(n12515) );
  XNOR2_X1 U14829 ( .A(n12515), .B(n12969), .ZN(n12594) );
  NAND2_X1 U14830 ( .A1(n12515), .A2(n12969), .ZN(n12516) );
  XNOR2_X1 U14831 ( .A(n12614), .B(n14769), .ZN(n12629) );
  INV_X1 U14832 ( .A(n12629), .ZN(n12518) );
  XNOR2_X1 U14833 ( .A(n12614), .B(n12634), .ZN(n12631) );
  NOR2_X1 U14834 ( .A1(n12631), .A2(n14775), .ZN(n12519) );
  INV_X1 U14835 ( .A(n12519), .ZN(n12517) );
  OAI21_X1 U14836 ( .B1(n12518), .B2(n12700), .A(n12517), .ZN(n12522) );
  NOR3_X1 U14837 ( .A1(n12519), .A2(n12968), .A3(n12629), .ZN(n12520) );
  AOI21_X1 U14838 ( .B1(n14775), .B2(n12631), .A(n12520), .ZN(n12521) );
  XNOR2_X1 U14839 ( .A(n14755), .B(n12614), .ZN(n12681) );
  NOR2_X1 U14840 ( .A1(n12681), .A2(n13262), .ZN(n12524) );
  NAND2_X1 U14841 ( .A1(n12681), .A2(n13262), .ZN(n12523) );
  XNOR2_X1 U14842 ( .A(n12579), .B(n12614), .ZN(n12525) );
  XNOR2_X1 U14843 ( .A(n12525), .B(n14759), .ZN(n12573) );
  XNOR2_X1 U14844 ( .A(n12736), .B(n12614), .ZN(n12527) );
  NAND2_X1 U14845 ( .A1(n12527), .A2(n13235), .ZN(n12725) );
  INV_X1 U14846 ( .A(n12527), .ZN(n12528) );
  NAND2_X1 U14847 ( .A1(n12528), .A2(n13263), .ZN(n12726) );
  INV_X1 U14848 ( .A(n12650), .ZN(n12531) );
  XOR2_X1 U14849 ( .A(n12614), .B(n13239), .Z(n12648) );
  INV_X1 U14850 ( .A(n12648), .ZN(n12530) );
  XNOR2_X1 U14851 ( .A(n13322), .B(n12614), .ZN(n12532) );
  XOR2_X1 U14852 ( .A(n12966), .B(n12532), .Z(n12657) );
  INV_X1 U14853 ( .A(n12532), .ZN(n12533) );
  NOR2_X1 U14854 ( .A1(n12533), .A2(n13234), .ZN(n12534) );
  AOI21_X2 U14855 ( .B1(n12658), .B2(n12657), .A(n12534), .ZN(n12709) );
  XNOR2_X1 U14856 ( .A(n12535), .B(n12548), .ZN(n12707) );
  NAND2_X1 U14857 ( .A1(n12707), .A2(n13222), .ZN(n12599) );
  XNOR2_X1 U14858 ( .A(n13309), .B(n12614), .ZN(n12540) );
  NAND2_X1 U14859 ( .A1(n12540), .A2(n13184), .ZN(n12537) );
  AND2_X1 U14860 ( .A1(n12599), .A2(n12537), .ZN(n12536) );
  XNOR2_X1 U14861 ( .A(n13305), .B(n12614), .ZN(n12544) );
  XNOR2_X1 U14862 ( .A(n12544), .B(n13200), .ZN(n12675) );
  INV_X1 U14863 ( .A(n12537), .ZN(n12542) );
  INV_X1 U14864 ( .A(n12707), .ZN(n12539) );
  NAND2_X1 U14865 ( .A1(n12539), .A2(n12538), .ZN(n12600) );
  XNOR2_X1 U14866 ( .A(n12540), .B(n13184), .ZN(n12601) );
  INV_X1 U14867 ( .A(n12601), .ZN(n12541) );
  AND2_X1 U14868 ( .A1(n12600), .A2(n12541), .ZN(n12603) );
  OR2_X1 U14869 ( .A1(n12542), .A2(n12603), .ZN(n12671) );
  AND2_X1 U14870 ( .A1(n12675), .A2(n12671), .ZN(n12543) );
  INV_X1 U14871 ( .A(n12544), .ZN(n12545) );
  NAND2_X1 U14872 ( .A1(n12545), .A2(n13200), .ZN(n12546) );
  XNOR2_X1 U14873 ( .A(n12872), .B(n12614), .ZN(n12547) );
  XOR2_X1 U14874 ( .A(n13185), .B(n12547), .Z(n12623) );
  XNOR2_X1 U14875 ( .A(n12695), .B(n12548), .ZN(n12549) );
  INV_X1 U14876 ( .A(n12550), .ZN(n12551) );
  XNOR2_X1 U14877 ( .A(n13155), .B(n12614), .ZN(n12553) );
  XNOR2_X1 U14878 ( .A(n12555), .B(n12553), .ZN(n12582) );
  NAND2_X1 U14879 ( .A1(n12582), .A2(n13164), .ZN(n12557) );
  INV_X1 U14880 ( .A(n12553), .ZN(n12554) );
  OR2_X1 U14881 ( .A1(n12555), .A2(n12554), .ZN(n12556) );
  NAND2_X1 U14882 ( .A1(n12557), .A2(n12556), .ZN(n12664) );
  XNOR2_X1 U14883 ( .A(n13289), .B(n12614), .ZN(n12558) );
  XOR2_X1 U14884 ( .A(n13151), .B(n12558), .Z(n12665) );
  NAND2_X1 U14885 ( .A1(n12664), .A2(n12665), .ZN(n12561) );
  INV_X1 U14886 ( .A(n12558), .ZN(n12559) );
  NAND2_X1 U14887 ( .A1(n12559), .A2(n12644), .ZN(n12560) );
  XNOR2_X1 U14888 ( .A(n13128), .B(n12614), .ZN(n12562) );
  XNOR2_X1 U14889 ( .A(n12562), .B(n13135), .ZN(n12641) );
  NAND2_X1 U14890 ( .A1(n12562), .A2(n13110), .ZN(n12563) );
  XNOR2_X1 U14891 ( .A(n12564), .B(n12614), .ZN(n12566) );
  XNOR2_X1 U14892 ( .A(n12566), .B(n13125), .ZN(n12716) );
  XNOR2_X1 U14893 ( .A(n12899), .B(n12614), .ZN(n12611) );
  XNOR2_X1 U14894 ( .A(n12611), .B(n12897), .ZN(n12612) );
  XNOR2_X1 U14895 ( .A(n12613), .B(n12612), .ZN(n12567) );
  NAND2_X1 U14896 ( .A1(n12567), .A2(n12673), .ZN(n12572) );
  AOI22_X1 U14897 ( .A1(n12731), .A2(n13125), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12568) );
  OAI21_X1 U14898 ( .B1(n12569), .B2(n12734), .A(n12568), .ZN(n12570) );
  AOI21_X1 U14899 ( .B1(n13099), .B2(n12729), .A(n12570), .ZN(n12571) );
  OAI211_X1 U14900 ( .C1(n13101), .C2(n12720), .A(n12572), .B(n12571), .ZN(
        P3_U3154) );
  XNOR2_X1 U14901 ( .A(n6690), .B(n12573), .ZN(n12581) );
  NAND2_X1 U14902 ( .A1(n12729), .A2(n13267), .ZN(n12577) );
  AOI21_X1 U14903 ( .B1(n12717), .B2(n13263), .A(n12575), .ZN(n12576) );
  OAI211_X1 U14904 ( .C1(n6878), .C2(n12719), .A(n12577), .B(n12576), .ZN(
        n12578) );
  AOI21_X1 U14905 ( .B1(n12737), .B2(n12579), .A(n12578), .ZN(n12580) );
  OAI21_X1 U14906 ( .B1(n12581), .B2(n12739), .A(n12580), .ZN(P3_U3155) );
  XNOR2_X1 U14907 ( .A(n12582), .B(n13136), .ZN(n12587) );
  NAND2_X1 U14908 ( .A1(n12729), .A2(n13156), .ZN(n12584) );
  AOI22_X1 U14909 ( .A1(n12717), .A2(n13151), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12583) );
  OAI211_X1 U14910 ( .C1(n13175), .C2(n12719), .A(n12584), .B(n12583), .ZN(
        n12585) );
  AOI21_X1 U14911 ( .B1(n13155), .B2(n12737), .A(n12585), .ZN(n12586) );
  OAI21_X1 U14912 ( .B1(n12587), .B2(n12739), .A(n12586), .ZN(P3_U3156) );
  AOI22_X1 U14913 ( .A1(n12737), .A2(n12588), .B1(n12731), .B2(n12970), .ZN(
        n12590) );
  OAI211_X1 U14914 ( .C1(n12700), .C2(n12734), .A(n12590), .B(n12589), .ZN(
        n12596) );
  INV_X1 U14915 ( .A(n12591), .ZN(n12592) );
  AOI211_X1 U14916 ( .C1(n12594), .C2(n12593), .A(n12739), .B(n12592), .ZN(
        n12595) );
  AOI211_X1 U14917 ( .C1(n12597), .C2(n12729), .A(n12596), .B(n12595), .ZN(
        n12598) );
  INV_X1 U14918 ( .A(n12598), .ZN(P3_U3157) );
  NAND2_X1 U14919 ( .A1(n12709), .A2(n12599), .ZN(n12604) );
  NAND2_X1 U14920 ( .A1(n12604), .A2(n12600), .ZN(n12602) );
  AOI21_X1 U14921 ( .B1(n12602), .B2(n12601), .A(n12739), .ZN(n12606) );
  NAND2_X1 U14922 ( .A1(n12604), .A2(n12603), .ZN(n12605) );
  NAND2_X1 U14923 ( .A1(n12606), .A2(n12605), .ZN(n12610) );
  NAND2_X1 U14924 ( .A1(n12731), .A2(n13222), .ZN(n12607) );
  NAND2_X1 U14925 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13068)
         );
  OAI211_X1 U14926 ( .C1(n13174), .C2(n12734), .A(n12607), .B(n13068), .ZN(
        n12608) );
  AOI21_X1 U14927 ( .B1(n12729), .B2(n13203), .A(n12608), .ZN(n12609) );
  OAI211_X1 U14928 ( .C1(n12720), .C2(n13309), .A(n12610), .B(n12609), .ZN(
        P3_U3159) );
  AOI22_X1 U14929 ( .A1(n12613), .A2(n12612), .B1(n13111), .B2(n12611), .ZN(
        n12616) );
  XOR2_X1 U14930 ( .A(n12614), .B(n12909), .Z(n12615) );
  XNOR2_X1 U14931 ( .A(n12616), .B(n12615), .ZN(n12621) );
  AOI22_X1 U14932 ( .A1(n12731), .A2(n12897), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12617) );
  OAI21_X1 U14933 ( .B1(n13089), .B2(n12734), .A(n12617), .ZN(n12619) );
  NOR2_X1 U14934 ( .A1(n13095), .A2(n12720), .ZN(n12618) );
  AOI211_X1 U14935 ( .C1(n13093), .C2(n12729), .A(n12619), .B(n12618), .ZN(
        n12620) );
  OAI21_X1 U14936 ( .B1(n12621), .B2(n12739), .A(n12620), .ZN(P3_U3160) );
  AOI21_X1 U14937 ( .B1(n12623), .B2(n12622), .A(n6488), .ZN(n12628) );
  NAND2_X1 U14938 ( .A1(n12729), .A2(n13178), .ZN(n12625) );
  AOI22_X1 U14939 ( .A1(n12731), .A2(n13200), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12624) );
  OAI211_X1 U14940 ( .C1(n13175), .C2(n12734), .A(n12625), .B(n12624), .ZN(
        n12626) );
  AOI21_X1 U14941 ( .B1(n12872), .B2(n12737), .A(n12626), .ZN(n12627) );
  OAI21_X1 U14942 ( .B1(n12628), .B2(n12739), .A(n12627), .ZN(P3_U3163) );
  XNOR2_X1 U14943 ( .A(n12630), .B(n12629), .ZN(n12699) );
  NOR2_X1 U14944 ( .A1(n12699), .A2(n12700), .ZN(n12698) );
  AOI21_X1 U14945 ( .B1(n12630), .B2(n12629), .A(n12698), .ZN(n12633) );
  XNOR2_X1 U14946 ( .A(n12631), .B(n14775), .ZN(n12632) );
  XNOR2_X1 U14947 ( .A(n12633), .B(n12632), .ZN(n12639) );
  AOI22_X1 U14948 ( .A1(n12737), .A2(n12634), .B1(n12731), .B2(n12968), .ZN(
        n12635) );
  NAND2_X1 U14949 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n12984)
         );
  OAI211_X1 U14950 ( .C1(n6878), .C2(n12734), .A(n12635), .B(n12984), .ZN(
        n12636) );
  AOI21_X1 U14951 ( .B1(n12637), .B2(n12729), .A(n12636), .ZN(n12638) );
  OAI21_X1 U14952 ( .B1(n12639), .B2(n12739), .A(n12638), .ZN(P3_U3164) );
  XOR2_X1 U14953 ( .A(n12641), .B(n12640), .Z(n12647) );
  NAND2_X1 U14954 ( .A1(n12729), .A2(n13129), .ZN(n12643) );
  AOI22_X1 U14955 ( .A1(n12717), .A2(n13125), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12642) );
  OAI211_X1 U14956 ( .C1(n12644), .C2(n12719), .A(n12643), .B(n12642), .ZN(
        n12645) );
  AOI21_X1 U14957 ( .B1(n13128), .B2(n12737), .A(n12645), .ZN(n12646) );
  OAI21_X1 U14958 ( .B1(n12647), .B2(n12739), .A(n12646), .ZN(P3_U3165) );
  XNOR2_X1 U14959 ( .A(n12648), .B(n13248), .ZN(n12649) );
  XNOR2_X1 U14960 ( .A(n12650), .B(n12649), .ZN(n12656) );
  NAND2_X1 U14961 ( .A1(n12729), .A2(n13240), .ZN(n12653) );
  NOR2_X1 U14962 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12651), .ZN(n13005) );
  AOI21_X1 U14963 ( .B1(n12717), .B2(n12966), .A(n13005), .ZN(n12652) );
  OAI211_X1 U14964 ( .C1(n13235), .C2(n12719), .A(n12653), .B(n12652), .ZN(
        n12654) );
  AOI21_X1 U14965 ( .B1(n12737), .B2(n13239), .A(n12654), .ZN(n12655) );
  OAI21_X1 U14966 ( .B1(n12656), .B2(n12739), .A(n12655), .ZN(P3_U3166) );
  XNOR2_X1 U14967 ( .A(n12658), .B(n12657), .ZN(n12663) );
  AND2_X1 U14968 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13025) );
  AOI21_X1 U14969 ( .B1(n12717), .B2(n13222), .A(n13025), .ZN(n12659) );
  OAI21_X1 U14970 ( .B1(n13248), .B2(n12719), .A(n12659), .ZN(n12661) );
  NOR2_X1 U14971 ( .A1(n13322), .A2(n12720), .ZN(n12660) );
  AOI211_X1 U14972 ( .C1(n13227), .C2(n12729), .A(n12661), .B(n12660), .ZN(
        n12662) );
  OAI21_X1 U14973 ( .B1(n12663), .B2(n12739), .A(n12662), .ZN(P3_U3168) );
  XOR2_X1 U14974 ( .A(n12665), .B(n12664), .Z(n12670) );
  AOI22_X1 U14975 ( .A1(n12717), .A2(n13135), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12666) );
  OAI21_X1 U14976 ( .B1(n13164), .B2(n12719), .A(n12666), .ZN(n12668) );
  NOR2_X1 U14977 ( .A1(n13289), .A2(n12720), .ZN(n12667) );
  AOI211_X1 U14978 ( .C1(n13141), .C2(n12729), .A(n12668), .B(n12667), .ZN(
        n12669) );
  OAI21_X1 U14979 ( .B1(n12670), .B2(n12739), .A(n12669), .ZN(P3_U3169) );
  INV_X1 U14980 ( .A(n13305), .ZN(n13192) );
  AND2_X1 U14981 ( .A1(n12672), .A2(n12671), .ZN(n12676) );
  OAI211_X1 U14982 ( .C1(n12676), .C2(n12675), .A(n12674), .B(n12673), .ZN(
        n12680) );
  AOI22_X1 U14983 ( .A1(n12717), .A2(n13185), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12677) );
  OAI21_X1 U14984 ( .B1(n13211), .B2(n12719), .A(n12677), .ZN(n12678) );
  AOI21_X1 U14985 ( .B1(n13190), .B2(n12729), .A(n12678), .ZN(n12679) );
  OAI211_X1 U14986 ( .C1(n13192), .C2(n12720), .A(n12680), .B(n12679), .ZN(
        P3_U3173) );
  XNOR2_X1 U14987 ( .A(n12681), .B(n13262), .ZN(n12682) );
  XNOR2_X1 U14988 ( .A(n12683), .B(n12682), .ZN(n12690) );
  NAND2_X1 U14989 ( .A1(n12729), .A2(n12684), .ZN(n12687) );
  AOI21_X1 U14990 ( .B1(n12717), .B2(n14759), .A(n12685), .ZN(n12686) );
  OAI211_X1 U14991 ( .C1(n14775), .C2(n12719), .A(n12687), .B(n12686), .ZN(
        n12688) );
  AOI21_X1 U14992 ( .B1(n13257), .B2(n12737), .A(n12688), .ZN(n12689) );
  OAI21_X1 U14993 ( .B1(n12690), .B2(n12739), .A(n12689), .ZN(P3_U3174) );
  XNOR2_X1 U14994 ( .A(n12691), .B(n6887), .ZN(n12697) );
  NAND2_X1 U14995 ( .A1(n12729), .A2(n13167), .ZN(n12693) );
  AOI22_X1 U14996 ( .A1(n12731), .A2(n13185), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12692) );
  OAI211_X1 U14997 ( .C1(n13164), .C2(n12734), .A(n12693), .B(n12692), .ZN(
        n12694) );
  AOI21_X1 U14998 ( .B1(n12695), .B2(n12737), .A(n12694), .ZN(n12696) );
  OAI21_X1 U14999 ( .B1(n12697), .B2(n12739), .A(n12696), .ZN(P3_U3175) );
  AOI211_X1 U15000 ( .C1(n12700), .C2(n12699), .A(n12739), .B(n12698), .ZN(
        n12701) );
  INV_X1 U15001 ( .A(n12701), .ZN(n12705) );
  INV_X1 U15002 ( .A(n14775), .ZN(n12967) );
  OAI22_X1 U15003 ( .A1(n12720), .A2(n14769), .B1(n14777), .B2(n12719), .ZN(
        n12702) );
  AOI211_X1 U15004 ( .C1(n12717), .C2(n12967), .A(n12703), .B(n12702), .ZN(
        n12704) );
  OAI211_X1 U15005 ( .C1(n14783), .C2(n12706), .A(n12705), .B(n12704), .ZN(
        P3_U3176) );
  XNOR2_X1 U15006 ( .A(n12707), .B(n13222), .ZN(n12708) );
  XNOR2_X1 U15007 ( .A(n12709), .B(n12708), .ZN(n12714) );
  NAND2_X1 U15008 ( .A1(n12731), .A2(n12966), .ZN(n12710) );
  NAND2_X1 U15009 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13048)
         );
  OAI211_X1 U15010 ( .C1(n13211), .C2(n12734), .A(n12710), .B(n13048), .ZN(
        n12712) );
  NOR2_X1 U15011 ( .A1(n13371), .A2(n12720), .ZN(n12711) );
  AOI211_X1 U15012 ( .C1(n13215), .C2(n12729), .A(n12712), .B(n12711), .ZN(
        n12713) );
  OAI21_X1 U15013 ( .B1(n12714), .B2(n12739), .A(n12713), .ZN(P3_U3178) );
  XOR2_X1 U15014 ( .A(n12716), .B(n12715), .Z(n12724) );
  AOI22_X1 U15015 ( .A1(n12717), .A2(n12897), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12718) );
  OAI21_X1 U15016 ( .B1(n13110), .B2(n12719), .A(n12718), .ZN(n12722) );
  NOR2_X1 U15017 ( .A1(n13348), .A2(n12720), .ZN(n12721) );
  AOI211_X1 U15018 ( .C1(n13117), .C2(n12729), .A(n12722), .B(n12721), .ZN(
        n12723) );
  OAI21_X1 U15019 ( .B1(n12724), .B2(n12739), .A(n12723), .ZN(P3_U3180) );
  NAND2_X1 U15020 ( .A1(n12726), .A2(n12725), .ZN(n12728) );
  XOR2_X1 U15021 ( .A(n12728), .B(n12727), .Z(n12740) );
  NAND2_X1 U15022 ( .A1(n12729), .A2(n13251), .ZN(n12733) );
  AOI21_X1 U15023 ( .B1(n12731), .B2(n14759), .A(n12730), .ZN(n12732) );
  OAI211_X1 U15024 ( .C1(n13248), .C2(n12734), .A(n12733), .B(n12732), .ZN(
        n12735) );
  AOI21_X1 U15025 ( .B1(n12737), .B2(n12736), .A(n12735), .ZN(n12738) );
  OAI21_X1 U15026 ( .B1(n12740), .B2(n12739), .A(n12738), .ZN(P3_U3181) );
  XNOR2_X1 U15027 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12745) );
  INV_X1 U15028 ( .A(SI_31_), .ZN(n13390) );
  OR2_X1 U15029 ( .A1(n6422), .A2(n13390), .ZN(n12746) );
  NAND2_X1 U15030 ( .A1(n12747), .A2(n12746), .ZN(n12756) );
  NAND2_X1 U15031 ( .A1(n12749), .A2(n12748), .ZN(n12752) );
  OR2_X1 U15032 ( .A1(n6422), .A2(n12750), .ZN(n12751) );
  AOI21_X1 U15033 ( .B1(n13339), .B2(n13081), .A(n12920), .ZN(n12753) );
  NAND2_X1 U15034 ( .A1(n13339), .A2(n12755), .ZN(n12912) );
  AND2_X1 U15035 ( .A1(n12918), .A2(n7405), .ZN(n12754) );
  OR2_X1 U15036 ( .A1(n13339), .A2(n12755), .ZN(n12925) );
  NOR2_X1 U15037 ( .A1(n13337), .A2(n12925), .ZN(n12757) );
  NAND2_X1 U15038 ( .A1(n12759), .A2(n12758), .ZN(n12760) );
  INV_X1 U15039 ( .A(n12762), .ZN(n12957) );
  INV_X1 U15040 ( .A(n12763), .ZN(n12764) );
  AOI22_X1 U15041 ( .A1(n12766), .A2(n12764), .B1(n13289), .B2(n13151), .ZN(
        n12765) );
  MUX2_X1 U15042 ( .A(n12766), .B(n12765), .S(n12919), .Z(n12888) );
  INV_X1 U15043 ( .A(n13140), .ZN(n12886) );
  INV_X1 U15044 ( .A(n12775), .ZN(n12767) );
  AOI21_X1 U15045 ( .B1(n15189), .B2(n12768), .A(n12767), .ZN(n12769) );
  MUX2_X1 U15046 ( .A(n12770), .B(n12769), .S(n12917), .Z(n12783) );
  NAND3_X1 U15047 ( .A1(n15193), .A2(n12771), .A3(n12962), .ZN(n12772) );
  OAI21_X1 U15048 ( .B1(n15190), .B2(n12773), .A(n12772), .ZN(n12776) );
  AOI21_X1 U15049 ( .B1(n12776), .B2(n12775), .A(n12774), .ZN(n12782) );
  NAND2_X1 U15050 ( .A1(n12785), .A2(n12777), .ZN(n12780) );
  NAND2_X1 U15051 ( .A1(n12784), .A2(n12778), .ZN(n12779) );
  MUX2_X1 U15052 ( .A(n12780), .B(n12779), .S(n12917), .Z(n12781) );
  AOI21_X1 U15053 ( .B1(n12783), .B2(n12782), .A(n12781), .ZN(n12792) );
  MUX2_X1 U15054 ( .A(n12785), .B(n12784), .S(n12919), .Z(n12786) );
  NAND2_X1 U15055 ( .A1(n12786), .A2(n12937), .ZN(n12791) );
  NAND2_X1 U15056 ( .A1(n12975), .A2(n12787), .ZN(n12788) );
  MUX2_X1 U15057 ( .A(n12789), .B(n12788), .S(n12917), .Z(n12790) );
  OAI211_X1 U15058 ( .C1(n12792), .C2(n12791), .A(n12931), .B(n12790), .ZN(
        n12797) );
  NAND2_X1 U15059 ( .A1(n12800), .A2(n12793), .ZN(n12794) );
  NAND2_X1 U15060 ( .A1(n12794), .A2(n12917), .ZN(n12796) );
  INV_X1 U15061 ( .A(n12799), .ZN(n12795) );
  AOI21_X1 U15062 ( .B1(n12797), .B2(n12796), .A(n12795), .ZN(n12804) );
  AOI21_X1 U15063 ( .B1(n12799), .B2(n12798), .A(n12917), .ZN(n12803) );
  INV_X1 U15064 ( .A(n12800), .ZN(n12801) );
  AOI21_X1 U15065 ( .B1(n12801), .B2(n12919), .A(n12933), .ZN(n12802) );
  OAI21_X1 U15066 ( .B1(n12804), .B2(n12803), .A(n12802), .ZN(n12810) );
  NAND2_X1 U15067 ( .A1(n12805), .A2(n12917), .ZN(n12808) );
  NAND2_X1 U15068 ( .A1(n12972), .A2(n12919), .ZN(n12807) );
  MUX2_X1 U15069 ( .A(n12808), .B(n12807), .S(n12806), .Z(n12809) );
  NAND3_X1 U15070 ( .A1(n12810), .A2(n12932), .A3(n12809), .ZN(n12814) );
  MUX2_X1 U15071 ( .A(n12812), .B(n12811), .S(n12917), .Z(n12813) );
  NAND4_X1 U15072 ( .A1(n12814), .A2(n12936), .A3(n12927), .A4(n12813), .ZN(
        n12826) );
  INV_X1 U15073 ( .A(n12815), .ZN(n12818) );
  INV_X1 U15074 ( .A(n12816), .ZN(n12817) );
  MUX2_X1 U15075 ( .A(n12818), .B(n12817), .S(n12917), .Z(n12824) );
  INV_X1 U15076 ( .A(n12819), .ZN(n12822) );
  INV_X1 U15077 ( .A(n12820), .ZN(n12821) );
  MUX2_X1 U15078 ( .A(n12822), .B(n12821), .S(n12917), .Z(n12823) );
  AOI21_X1 U15079 ( .B1(n12927), .B2(n12824), .A(n12823), .ZN(n12825) );
  NAND4_X1 U15080 ( .A1(n12826), .A2(n8056), .A3(n12938), .A4(n12825), .ZN(
        n12836) );
  NAND2_X1 U15081 ( .A1(n12831), .A2(n12827), .ZN(n12828) );
  NAND2_X1 U15082 ( .A1(n12828), .A2(n12830), .ZN(n12834) );
  NAND2_X1 U15083 ( .A1(n12968), .A2(n14769), .ZN(n12829) );
  NAND2_X1 U15084 ( .A1(n12830), .A2(n12829), .ZN(n12832) );
  NAND2_X1 U15085 ( .A1(n12832), .A2(n12831), .ZN(n12833) );
  MUX2_X1 U15086 ( .A(n12834), .B(n12833), .S(n12917), .Z(n12835) );
  NAND3_X1 U15087 ( .A1(n12836), .A2(n14758), .A3(n12835), .ZN(n12842) );
  INV_X1 U15088 ( .A(n12837), .ZN(n12838) );
  MUX2_X1 U15089 ( .A(n12839), .B(n12838), .S(n12917), .Z(n12840) );
  NOR2_X1 U15090 ( .A1(n13260), .A2(n12840), .ZN(n12841) );
  NAND2_X1 U15091 ( .A1(n12842), .A2(n12841), .ZN(n12846) );
  INV_X1 U15092 ( .A(n13249), .ZN(n12942) );
  MUX2_X1 U15093 ( .A(n12844), .B(n12843), .S(n12919), .Z(n12845) );
  NAND3_X1 U15094 ( .A1(n12846), .A2(n12942), .A3(n12845), .ZN(n12851) );
  NAND2_X1 U15095 ( .A1(n12854), .A2(n12847), .ZN(n12848) );
  NAND2_X1 U15096 ( .A1(n12848), .A2(n12919), .ZN(n12850) );
  INV_X1 U15097 ( .A(n12853), .ZN(n12849) );
  AOI21_X1 U15098 ( .B1(n12851), .B2(n12850), .A(n12849), .ZN(n12856) );
  AOI21_X1 U15099 ( .B1(n12853), .B2(n12852), .A(n12919), .ZN(n12855) );
  OAI22_X1 U15100 ( .A1(n12856), .A2(n12855), .B1(n12919), .B2(n12854), .ZN(
        n12862) );
  INV_X1 U15101 ( .A(n12863), .ZN(n12861) );
  AND2_X1 U15102 ( .A1(n12858), .A2(n12917), .ZN(n12859) );
  OAI211_X1 U15103 ( .C1(n12861), .C2(n12860), .A(n12869), .B(n12859), .ZN(
        n12865) );
  AOI22_X1 U15104 ( .A1(n12862), .A2(n13225), .B1(n7048), .B2(n12865), .ZN(
        n12867) );
  NAND3_X1 U15105 ( .A1(n12868), .A2(n12919), .A3(n12863), .ZN(n12864) );
  NAND2_X1 U15106 ( .A1(n12865), .A2(n12864), .ZN(n12866) );
  OAI21_X1 U15107 ( .B1(n12867), .B2(n13214), .A(n12866), .ZN(n12871) );
  MUX2_X1 U15108 ( .A(n12869), .B(n12868), .S(n12917), .Z(n12870) );
  NAND3_X1 U15109 ( .A1(n12871), .A2(n13188), .A3(n12870), .ZN(n12876) );
  XNOR2_X1 U15110 ( .A(n12872), .B(n13185), .ZN(n13177) );
  MUX2_X1 U15111 ( .A(n12874), .B(n12873), .S(n12917), .Z(n12875) );
  NAND3_X1 U15112 ( .A1(n12876), .A2(n13177), .A3(n12875), .ZN(n12879) );
  MUX2_X1 U15113 ( .A(n6431), .B(n12877), .S(n12917), .Z(n12878) );
  NAND3_X1 U15114 ( .A1(n12879), .A2(n13165), .A3(n12878), .ZN(n12882) );
  MUX2_X1 U15115 ( .A(n6471), .B(n12880), .S(n12917), .Z(n12881) );
  NAND3_X1 U15116 ( .A1(n12882), .A2(n13148), .A3(n12881), .ZN(n12884) );
  NAND3_X1 U15117 ( .A1(n13155), .A2(n13164), .A3(n12917), .ZN(n12883) );
  NAND2_X1 U15118 ( .A1(n12884), .A2(n12883), .ZN(n12885) );
  NAND2_X1 U15119 ( .A1(n12886), .A2(n12885), .ZN(n12887) );
  NAND3_X1 U15120 ( .A1(n12888), .A2(n12926), .A3(n12887), .ZN(n12892) );
  MUX2_X1 U15121 ( .A(n12890), .B(n12889), .S(n12917), .Z(n12891) );
  NAND3_X1 U15122 ( .A1(n13109), .A2(n12892), .A3(n12891), .ZN(n12896) );
  MUX2_X1 U15123 ( .A(n12894), .B(n12893), .S(n12919), .Z(n12895) );
  NAND2_X1 U15124 ( .A1(n12896), .A2(n12895), .ZN(n12901) );
  NAND2_X1 U15125 ( .A1(n12897), .A2(n12919), .ZN(n12898) );
  NOR2_X1 U15126 ( .A1(n12899), .A2(n12898), .ZN(n12900) );
  AOI21_X1 U15127 ( .B1(n12947), .B2(n12901), .A(n12900), .ZN(n12910) );
  INV_X1 U15128 ( .A(n12902), .ZN(n12903) );
  NAND2_X1 U15129 ( .A1(n12904), .A2(n12903), .ZN(n12905) );
  NAND2_X1 U15130 ( .A1(n12905), .A2(n12907), .ZN(n12906) );
  MUX2_X1 U15131 ( .A(n12907), .B(n12906), .S(n12917), .Z(n12908) );
  OAI21_X1 U15132 ( .B1(n12910), .B2(n12909), .A(n12908), .ZN(n12911) );
  NAND2_X1 U15133 ( .A1(n12911), .A2(n12949), .ZN(n12913) );
  NAND3_X1 U15134 ( .A1(n12913), .A2(n12912), .A3(n12925), .ZN(n12921) );
  INV_X1 U15135 ( .A(n12914), .ZN(n12915) );
  NOR2_X1 U15136 ( .A1(n12921), .A2(n12915), .ZN(n12916) );
  AOI211_X1 U15137 ( .C1(n12917), .C2(n12925), .A(n12952), .B(n12916), .ZN(
        n12924) );
  INV_X1 U15138 ( .A(n12918), .ZN(n12922) );
  NOR4_X1 U15139 ( .A1(n12922), .A2(n12921), .A3(n12920), .A4(n12919), .ZN(
        n12923) );
  NOR3_X1 U15140 ( .A1(n12924), .A2(n7404), .A3(n12923), .ZN(n12956) );
  INV_X1 U15141 ( .A(n12925), .ZN(n12951) );
  NAND4_X1 U15142 ( .A1(n12929), .A2(n12928), .A3(n15189), .A4(n12927), .ZN(
        n12935) );
  NAND4_X1 U15143 ( .A1(n12932), .A2(n15175), .A3(n12931), .A4(n12930), .ZN(
        n12934) );
  NOR3_X1 U15144 ( .A1(n12935), .A2(n12934), .A3(n12933), .ZN(n12939) );
  NAND4_X1 U15145 ( .A1(n12939), .A2(n12938), .A3(n12937), .A4(n12936), .ZN(
        n12940) );
  INV_X1 U15146 ( .A(n14758), .ZN(n14756) );
  NOR4_X1 U15147 ( .A1(n13260), .A2(n14772), .A3(n12940), .A4(n14756), .ZN(
        n12941) );
  NAND4_X1 U15148 ( .A1(n13237), .A2(n13225), .A3(n12942), .A4(n12941), .ZN(
        n12943) );
  NOR4_X1 U15149 ( .A1(n12944), .A2(n13214), .A3(n13198), .A4(n12943), .ZN(
        n12945) );
  NAND4_X1 U15150 ( .A1(n13148), .A2(n13165), .A3(n12945), .A4(n13177), .ZN(
        n12946) );
  NOR4_X1 U15151 ( .A1(n13106), .A2(n13124), .A3(n13140), .A4(n12946), .ZN(
        n12948) );
  NAND4_X1 U15152 ( .A1(n12949), .A2(n13087), .A3(n12948), .A4(n12947), .ZN(
        n12950) );
  OAI22_X1 U15153 ( .A1(n12956), .A2(n15200), .B1(n12954), .B2(n12953), .ZN(
        n12955) );
  AOI21_X1 U15154 ( .B1(n12957), .B2(n12956), .A(n12955), .ZN(n12958) );
  INV_X1 U15155 ( .A(n12959), .ZN(n12963) );
  INV_X1 U15156 ( .A(P3_B_REG_SCAN_IN), .ZN(n13742) );
  NOR2_X1 U15157 ( .A1(n12960), .A2(n13056), .ZN(n12961) );
  AOI211_X1 U15158 ( .C1(n12963), .C2(n12962), .A(n13742), .B(n12961), .ZN(
        n12964) );
  MUX2_X1 U15159 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12965), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15160 ( .A(n13125), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12976), .Z(
        P3_U3517) );
  MUX2_X1 U15161 ( .A(n13135), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12976), .Z(
        P3_U3516) );
  MUX2_X1 U15162 ( .A(n13151), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12976), .Z(
        P3_U3515) );
  MUX2_X1 U15163 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n13136), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U15164 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n6887), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15165 ( .A(n13185), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12976), .Z(
        P3_U3512) );
  MUX2_X1 U15166 ( .A(n13200), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12976), .Z(
        P3_U3511) );
  MUX2_X1 U15167 ( .A(n13184), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12976), .Z(
        P3_U3510) );
  MUX2_X1 U15168 ( .A(n13222), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12976), .Z(
        P3_U3509) );
  MUX2_X1 U15169 ( .A(n12966), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12976), .Z(
        P3_U3508) );
  MUX2_X1 U15170 ( .A(n13221), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12976), .Z(
        P3_U3507) );
  MUX2_X1 U15171 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n13263), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U15172 ( .A(n14759), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12976), .Z(
        P3_U3505) );
  MUX2_X1 U15173 ( .A(n13262), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12976), .Z(
        P3_U3504) );
  MUX2_X1 U15174 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12967), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15175 ( .A(n12968), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12976), .Z(
        P3_U3502) );
  MUX2_X1 U15176 ( .A(n12969), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12976), .Z(
        P3_U3501) );
  MUX2_X1 U15177 ( .A(n12970), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12976), .Z(
        P3_U3500) );
  MUX2_X1 U15178 ( .A(n12971), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12976), .Z(
        P3_U3499) );
  MUX2_X1 U15179 ( .A(n12972), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12976), .Z(
        P3_U3498) );
  MUX2_X1 U15180 ( .A(n12973), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12976), .Z(
        P3_U3497) );
  MUX2_X1 U15181 ( .A(n12974), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12976), .Z(
        P3_U3496) );
  MUX2_X1 U15182 ( .A(n12975), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12976), .Z(
        P3_U3495) );
  MUX2_X1 U15183 ( .A(n15194), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12976), .Z(
        P3_U3493) );
  MUX2_X1 U15184 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n15173), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15185 ( .A(n15193), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12976), .Z(
        P3_U3491) );
  OAI211_X1 U15186 ( .C1(n12979), .C2(n12978), .A(n12977), .B(n15146), .ZN(
        n12994) );
  OAI21_X1 U15187 ( .B1(n12982), .B2(n12981), .A(n12980), .ZN(n12987) );
  NAND2_X1 U15188 ( .A1(n15113), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n12983) );
  OAI211_X1 U15189 ( .C1(n15150), .C2(n12985), .A(n12984), .B(n12983), .ZN(
        n12986) );
  AOI21_X1 U15190 ( .B1(n12987), .B2(n13023), .A(n12986), .ZN(n12993) );
  OAI21_X1 U15191 ( .B1(n12990), .B2(n12989), .A(n12988), .ZN(n12991) );
  NAND2_X1 U15192 ( .A1(n12991), .A2(n15154), .ZN(n12992) );
  NAND3_X1 U15193 ( .A1(n12994), .A2(n12993), .A3(n12992), .ZN(P3_U3194) );
  NAND2_X1 U15194 ( .A1(n13010), .A2(n12995), .ZN(n12997) );
  NAND2_X1 U15195 ( .A1(n12997), .A2(n12996), .ZN(n13000) );
  INV_X1 U15196 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12998) );
  MUX2_X1 U15197 ( .A(n12998), .B(P3_REG2_REG_16__SCAN_IN), .S(n13018), .Z(
        n12999) );
  NAND2_X1 U15198 ( .A1(n13000), .A2(n12999), .ZN(n13017) );
  OAI21_X1 U15199 ( .B1(n13000), .B2(n12999), .A(n13017), .ZN(n13015) );
  XNOR2_X1 U15200 ( .A(n13018), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n13020) );
  NAND2_X1 U15201 ( .A1(n13010), .A2(n13001), .ZN(n13003) );
  NAND2_X1 U15202 ( .A1(n13003), .A2(n13002), .ZN(n13021) );
  XOR2_X1 U15203 ( .A(n13020), .B(n13021), .Z(n13007) );
  NOR2_X1 U15204 ( .A1(n15150), .A2(n13029), .ZN(n13004) );
  AOI211_X1 U15205 ( .C1(n15113), .C2(P3_ADDR_REG_16__SCAN_IN), .A(n13005), 
        .B(n13004), .ZN(n13006) );
  OAI21_X1 U15206 ( .B1(n13007), .B2(n15140), .A(n13006), .ZN(n13014) );
  MUX2_X1 U15207 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n13037), .Z(n13030) );
  XOR2_X1 U15208 ( .A(n13018), .B(n13030), .Z(n13011) );
  AOI211_X1 U15209 ( .C1(n13012), .C2(n13011), .A(n13078), .B(n13028), .ZN(
        n13013) );
  AOI211_X1 U15210 ( .C1(n15154), .C2(n13015), .A(n13014), .B(n13013), .ZN(
        n13016) );
  INV_X1 U15211 ( .A(n13016), .ZN(P3_U3198) );
  OAI21_X1 U15212 ( .B1(n13018), .B2(n12998), .A(n13017), .ZN(n13043) );
  OAI21_X1 U15213 ( .B1(P3_REG2_REG_17__SCAN_IN), .B2(n13019), .A(n13042), 
        .ZN(n13035) );
  XNOR2_X1 U15214 ( .A(n13046), .B(n13044), .ZN(n13022) );
  NAND2_X1 U15215 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n13022), .ZN(n13045) );
  OAI21_X1 U15216 ( .B1(n13022), .B2(P3_REG1_REG_17__SCAN_IN), .A(n13045), 
        .ZN(n13024) );
  NAND2_X1 U15217 ( .A1(n13024), .A2(n13023), .ZN(n13027) );
  AOI21_X1 U15218 ( .B1(n15113), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n13025), 
        .ZN(n13026) );
  OAI211_X1 U15219 ( .C1(n15150), .C2(n13044), .A(n13027), .B(n13026), .ZN(
        n13034) );
  AOI21_X1 U15220 ( .B1(n13030), .B2(n13029), .A(n13028), .ZN(n13032) );
  MUX2_X1 U15221 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13037), .Z(n13039) );
  XNOR2_X1 U15222 ( .A(n13039), .B(n13044), .ZN(n13031) );
  NOR2_X1 U15223 ( .A1(n13032), .A2(n13031), .ZN(n13038) );
  AOI211_X1 U15224 ( .C1(n13032), .C2(n13031), .A(n13078), .B(n13038), .ZN(
        n13033) );
  AOI211_X1 U15225 ( .C1(n13035), .C2(n15154), .A(n13034), .B(n13033), .ZN(
        n13036) );
  INV_X1 U15226 ( .A(n13036), .ZN(P3_U3199) );
  MUX2_X1 U15227 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13037), .Z(n13041) );
  NOR2_X1 U15228 ( .A1(n13040), .A2(n13041), .ZN(n13054) );
  AOI21_X1 U15229 ( .B1(n13041), .B2(n13040), .A(n13054), .ZN(n13053) );
  XOR2_X1 U15230 ( .A(P3_REG2_REG_18__SCAN_IN), .B(n13058), .Z(n13059) );
  XNOR2_X1 U15231 ( .A(n13060), .B(n13059), .ZN(n13051) );
  XNOR2_X1 U15232 ( .A(n13058), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n13064) );
  OAI21_X1 U15233 ( .B1(n13046), .B2(n6581), .A(n13045), .ZN(n13065) );
  NOR2_X1 U15234 ( .A1(n6468), .A2(n15140), .ZN(n13050) );
  NAND2_X1 U15235 ( .A1(n15113), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n13047) );
  OAI211_X1 U15236 ( .C1(n15150), .C2(n13063), .A(n13048), .B(n13047), .ZN(
        n13049) );
  AOI211_X1 U15237 ( .C1(n13051), .C2(n15154), .A(n13050), .B(n13049), .ZN(
        n13052) );
  OAI21_X1 U15238 ( .B1(n13053), .B2(n13078), .A(n13052), .ZN(P3_U3200) );
  XNOR2_X1 U15239 ( .A(n13072), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13066) );
  XNOR2_X1 U15240 ( .A(n13072), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13061) );
  MUX2_X1 U15241 ( .A(n13066), .B(n13061), .S(n13056), .Z(n13057) );
  INV_X1 U15242 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13686) );
  OAI22_X1 U15243 ( .A1(n13060), .A2(n13059), .B1(n13058), .B2(n13686), .ZN(
        n13062) );
  XNOR2_X1 U15244 ( .A(n13062), .B(n13061), .ZN(n13076) );
  AOI22_X1 U15245 ( .A1(n13065), .A2(n13064), .B1(P3_REG1_REG_18__SCAN_IN), 
        .B2(n13063), .ZN(n13067) );
  XNOR2_X1 U15246 ( .A(n13067), .B(n13066), .ZN(n13074) );
  OAI21_X1 U15247 ( .B1(n15157), .B2(n13069), .A(n13068), .ZN(n13070) );
  AOI21_X1 U15248 ( .B1(n13072), .B2(n13071), .A(n13070), .ZN(n13073) );
  OAI21_X1 U15249 ( .B1(n13074), .B2(n15140), .A(n13073), .ZN(n13075) );
  AOI21_X1 U15250 ( .B1(n13076), .B2(n15154), .A(n13075), .ZN(n13077) );
  OAI21_X1 U15251 ( .B1(n13079), .B2(n13078), .A(n13077), .ZN(P3_U3201) );
  AOI21_X1 U15252 ( .B1(n13082), .B2(n13335), .A(n15206), .ZN(n13084) );
  AOI21_X1 U15253 ( .B1(n15206), .B2(P3_REG2_REG_31__SCAN_IN), .A(n13084), 
        .ZN(n13083) );
  OAI21_X1 U15254 ( .B1(n13337), .B2(n15165), .A(n13083), .ZN(P3_U3202) );
  INV_X1 U15255 ( .A(n13339), .ZN(n13276) );
  AOI21_X1 U15256 ( .B1(n15206), .B2(P3_REG2_REG_30__SCAN_IN), .A(n13084), 
        .ZN(n13085) );
  OAI21_X1 U15257 ( .B1(n13276), .B2(n15165), .A(n13085), .ZN(P3_U3203) );
  XNOR2_X1 U15258 ( .A(n13086), .B(n13087), .ZN(n13280) );
  AOI21_X1 U15259 ( .B1(n13088), .B2(n13087), .A(n15198), .ZN(n13092) );
  OAI22_X1 U15260 ( .A1(n13111), .A2(n14778), .B1(n13089), .B2(n14776), .ZN(
        n13090) );
  AOI21_X1 U15261 ( .B1(n13092), .B2(n13091), .A(n13090), .ZN(n13279) );
  INV_X1 U15262 ( .A(n13279), .ZN(n13097) );
  AOI22_X1 U15263 ( .A1(n15206), .A2(P3_REG2_REG_28__SCAN_IN), .B1(n15201), 
        .B2(n13093), .ZN(n13094) );
  OAI21_X1 U15264 ( .B1(n13095), .B2(n15165), .A(n13094), .ZN(n13096) );
  AOI21_X1 U15265 ( .B1(n13097), .B2(n15204), .A(n13096), .ZN(n13098) );
  OAI21_X1 U15266 ( .B1(n13280), .B2(n13207), .A(n13098), .ZN(P3_U3205) );
  AOI22_X1 U15267 ( .A1(n15206), .A2(P3_REG2_REG_27__SCAN_IN), .B1(n15201), 
        .B2(n13099), .ZN(n13100) );
  OAI21_X1 U15268 ( .B1(n13101), .B2(n15165), .A(n13100), .ZN(n13102) );
  AOI21_X1 U15269 ( .B1(n13103), .B2(n15204), .A(n13102), .ZN(n13104) );
  OAI21_X1 U15270 ( .B1(n13105), .B2(n13207), .A(n13104), .ZN(P3_U3206) );
  XNOR2_X1 U15271 ( .A(n13107), .B(n13106), .ZN(n13115) );
  XNOR2_X1 U15272 ( .A(n13108), .B(n13109), .ZN(n13113) );
  OAI22_X1 U15273 ( .A1(n13111), .A2(n14776), .B1(n13110), .B2(n14778), .ZN(
        n13112) );
  AOI21_X1 U15274 ( .B1(n13113), .B2(n14762), .A(n13112), .ZN(n13114) );
  OAI21_X1 U15275 ( .B1(n15177), .B2(n13115), .A(n13114), .ZN(n13281) );
  INV_X1 U15276 ( .A(n13281), .ZN(n13121) );
  INV_X1 U15277 ( .A(n13115), .ZN(n13282) );
  INV_X1 U15278 ( .A(n13116), .ZN(n15202) );
  AOI22_X1 U15279 ( .A1(n15206), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n15201), 
        .B2(n13117), .ZN(n13118) );
  OAI21_X1 U15280 ( .B1(n13348), .B2(n15165), .A(n13118), .ZN(n13119) );
  AOI21_X1 U15281 ( .B1(n13282), .B2(n15202), .A(n13119), .ZN(n13120) );
  OAI21_X1 U15282 ( .B1(n13121), .B2(n15206), .A(n13120), .ZN(P3_U3207) );
  XNOR2_X1 U15283 ( .A(n13122), .B(n13124), .ZN(n13286) );
  INV_X1 U15284 ( .A(n13286), .ZN(n13133) );
  OAI211_X1 U15285 ( .C1(n6505), .C2(n13124), .A(n14762), .B(n13123), .ZN(
        n13127) );
  AOI22_X1 U15286 ( .A1(n15195), .A2(n13125), .B1(n13151), .B2(n15192), .ZN(
        n13126) );
  NAND2_X1 U15287 ( .A1(n13127), .A2(n13126), .ZN(n13285) );
  INV_X1 U15288 ( .A(n13128), .ZN(n13352) );
  AOI22_X1 U15289 ( .A1(n15206), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n15201), 
        .B2(n13129), .ZN(n13130) );
  OAI21_X1 U15290 ( .B1(n13352), .B2(n15165), .A(n13130), .ZN(n13131) );
  AOI21_X1 U15291 ( .B1(n13285), .B2(n15204), .A(n13131), .ZN(n13132) );
  OAI21_X1 U15292 ( .B1(n13207), .B2(n13133), .A(n13132), .ZN(P3_U3208) );
  XNOR2_X1 U15293 ( .A(n13134), .B(n13140), .ZN(n13137) );
  AOI222_X1 U15294 ( .A1(n14762), .A2(n13137), .B1(n13136), .B2(n15192), .C1(
        n13135), .C2(n15195), .ZN(n13292) );
  AOI21_X1 U15295 ( .B1(n13140), .B2(n13139), .A(n13138), .ZN(n13293) );
  INV_X1 U15296 ( .A(n13293), .ZN(n13144) );
  AOI22_X1 U15297 ( .A1(n15206), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15201), 
        .B2(n13141), .ZN(n13142) );
  OAI21_X1 U15298 ( .B1(n13289), .B2(n15165), .A(n13142), .ZN(n13143) );
  AOI21_X1 U15299 ( .B1(n13144), .B2(n13270), .A(n13143), .ZN(n13145) );
  OAI21_X1 U15300 ( .B1(n13292), .B2(n15206), .A(n13145), .ZN(P3_U3209) );
  OAI21_X1 U15301 ( .B1(n13147), .B2(n13148), .A(n13146), .ZN(n13154) );
  XNOR2_X1 U15302 ( .A(n13149), .B(n13148), .ZN(n13150) );
  NAND2_X1 U15303 ( .A1(n13150), .A2(n14762), .ZN(n13153) );
  AOI22_X1 U15304 ( .A1(n6887), .A2(n15192), .B1(n15195), .B2(n13151), .ZN(
        n13152) );
  OAI211_X1 U15305 ( .C1(n15177), .C2(n13154), .A(n13153), .B(n13152), .ZN(
        n13294) );
  INV_X1 U15306 ( .A(n13294), .ZN(n13160) );
  INV_X1 U15307 ( .A(n13154), .ZN(n13295) );
  INV_X1 U15308 ( .A(n13155), .ZN(n13357) );
  AOI22_X1 U15309 ( .A1(n15206), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15201), 
        .B2(n13156), .ZN(n13157) );
  OAI21_X1 U15310 ( .B1(n13357), .B2(n15165), .A(n13157), .ZN(n13158) );
  AOI21_X1 U15311 ( .B1(n13295), .B2(n15202), .A(n13158), .ZN(n13159) );
  OAI21_X1 U15312 ( .B1(n13160), .B2(n15206), .A(n13159), .ZN(P3_U3210) );
  XOR2_X1 U15313 ( .A(n13165), .B(n13161), .Z(n13162) );
  OAI222_X1 U15314 ( .A1(n14776), .A2(n13164), .B1(n14778), .B2(n13163), .C1(
        n13162), .C2(n15198), .ZN(n13297) );
  INV_X1 U15315 ( .A(n13297), .ZN(n13171) );
  XNOR2_X1 U15316 ( .A(n13166), .B(n13165), .ZN(n13298) );
  AOI22_X1 U15317 ( .A1(n15206), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15201), 
        .B2(n13167), .ZN(n13168) );
  OAI21_X1 U15318 ( .B1(n13361), .B2(n15165), .A(n13168), .ZN(n13169) );
  AOI21_X1 U15319 ( .B1(n13298), .B2(n13270), .A(n13169), .ZN(n13170) );
  OAI21_X1 U15320 ( .B1(n13171), .B2(n15206), .A(n13170), .ZN(P3_U3211) );
  XNOR2_X1 U15321 ( .A(n13172), .B(n13177), .ZN(n13173) );
  OAI222_X1 U15322 ( .A1(n14776), .A2(n13175), .B1(n14778), .B2(n13174), .C1(
        n15198), .C2(n13173), .ZN(n13301) );
  INV_X1 U15323 ( .A(n13301), .ZN(n13182) );
  XOR2_X1 U15324 ( .A(n13177), .B(n13176), .Z(n13302) );
  AOI22_X1 U15325 ( .A1(n15206), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15201), 
        .B2(n13178), .ZN(n13179) );
  OAI21_X1 U15326 ( .B1(n13365), .B2(n15165), .A(n13179), .ZN(n13180) );
  AOI21_X1 U15327 ( .B1(n13302), .B2(n13270), .A(n13180), .ZN(n13181) );
  OAI21_X1 U15328 ( .B1(n13182), .B2(n15206), .A(n13181), .ZN(P3_U3212) );
  XNOR2_X1 U15329 ( .A(n13183), .B(n13188), .ZN(n13186) );
  AOI222_X1 U15330 ( .A1(n14762), .A2(n13186), .B1(n13185), .B2(n15195), .C1(
        n13184), .C2(n15192), .ZN(n13307) );
  OAI21_X1 U15331 ( .B1(n13189), .B2(n13188), .A(n13187), .ZN(n13308) );
  INV_X1 U15332 ( .A(n13308), .ZN(n13194) );
  AOI22_X1 U15333 ( .A1(n15206), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15201), 
        .B2(n13190), .ZN(n13191) );
  OAI21_X1 U15334 ( .B1(n13192), .B2(n15165), .A(n13191), .ZN(n13193) );
  AOI21_X1 U15335 ( .B1(n13194), .B2(n13270), .A(n13193), .ZN(n13195) );
  OAI21_X1 U15336 ( .B1(n13307), .B2(n15206), .A(n13195), .ZN(P3_U3213) );
  XNOR2_X1 U15337 ( .A(n13196), .B(n13198), .ZN(n13314) );
  OAI211_X1 U15338 ( .C1(n13199), .C2(n13198), .A(n13197), .B(n14762), .ZN(
        n13202) );
  AOI22_X1 U15339 ( .A1(n15192), .A2(n13222), .B1(n13200), .B2(n15195), .ZN(
        n13201) );
  NAND2_X1 U15340 ( .A1(n13202), .A2(n13201), .ZN(n13310) );
  AOI22_X1 U15341 ( .A1(n15206), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15201), 
        .B2(n13203), .ZN(n13204) );
  OAI21_X1 U15342 ( .B1(n13309), .B2(n15165), .A(n13204), .ZN(n13205) );
  AOI21_X1 U15343 ( .B1(n13310), .B2(n15204), .A(n13205), .ZN(n13206) );
  OAI21_X1 U15344 ( .B1(n13314), .B2(n13207), .A(n13206), .ZN(P3_U3214) );
  AOI21_X1 U15345 ( .B1(n13209), .B2(n13208), .A(n6545), .ZN(n13210) );
  OAI222_X1 U15346 ( .A1(n14776), .A2(n13211), .B1(n14778), .B2(n13234), .C1(
        n15198), .C2(n13210), .ZN(n13315) );
  INV_X1 U15347 ( .A(n13315), .ZN(n13219) );
  AOI21_X1 U15348 ( .B1(n13214), .B2(n13213), .A(n13212), .ZN(n13316) );
  AOI22_X1 U15349 ( .A1(n15206), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15201), 
        .B2(n13215), .ZN(n13216) );
  OAI21_X1 U15350 ( .B1(n13371), .B2(n15165), .A(n13216), .ZN(n13217) );
  AOI21_X1 U15351 ( .B1(n13316), .B2(n13270), .A(n13217), .ZN(n13218) );
  OAI21_X1 U15352 ( .B1(n13219), .B2(n15206), .A(n13218), .ZN(P3_U3215) );
  XOR2_X1 U15353 ( .A(n13225), .B(n13220), .Z(n13223) );
  AOI222_X1 U15354 ( .A1(n14762), .A2(n13223), .B1(n13222), .B2(n15195), .C1(
        n13221), .C2(n15192), .ZN(n13321) );
  OAI21_X1 U15355 ( .B1(n13226), .B2(n13225), .A(n13224), .ZN(n13319) );
  AOI22_X1 U15356 ( .A1(n15206), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15201), 
        .B2(n13227), .ZN(n13228) );
  OAI21_X1 U15357 ( .B1(n13322), .B2(n15165), .A(n13228), .ZN(n13229) );
  AOI21_X1 U15358 ( .B1(n13319), .B2(n13270), .A(n13229), .ZN(n13230) );
  OAI21_X1 U15359 ( .B1(n13321), .B2(n15206), .A(n13230), .ZN(P3_U3216) );
  XNOR2_X1 U15360 ( .A(n13232), .B(n13231), .ZN(n13233) );
  OAI222_X1 U15361 ( .A1(n14778), .A2(n13235), .B1(n14776), .B2(n13234), .C1(
        n13233), .C2(n15198), .ZN(n13323) );
  INV_X1 U15362 ( .A(n13323), .ZN(n13244) );
  OAI21_X1 U15363 ( .B1(n13238), .B2(n13237), .A(n13236), .ZN(n13324) );
  INV_X1 U15364 ( .A(n13239), .ZN(n13376) );
  AOI22_X1 U15365 ( .A1(n15206), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15201), 
        .B2(n13240), .ZN(n13241) );
  OAI21_X1 U15366 ( .B1(n13376), .B2(n15165), .A(n13241), .ZN(n13242) );
  AOI21_X1 U15367 ( .B1(n13324), .B2(n13270), .A(n13242), .ZN(n13243) );
  OAI21_X1 U15368 ( .B1(n13244), .B2(n15206), .A(n13243), .ZN(P3_U3217) );
  XNOR2_X1 U15369 ( .A(n13245), .B(n13249), .ZN(n13246) );
  OAI222_X1 U15370 ( .A1(n14776), .A2(n13248), .B1(n14778), .B2(n13247), .C1(
        n13246), .C2(n15198), .ZN(n13326) );
  INV_X1 U15371 ( .A(n13326), .ZN(n13255) );
  XNOR2_X1 U15372 ( .A(n13250), .B(n13249), .ZN(n13327) );
  AOI22_X1 U15373 ( .A1(n15206), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15201), 
        .B2(n13251), .ZN(n13252) );
  OAI21_X1 U15374 ( .B1(n15165), .B2(n13380), .A(n13252), .ZN(n13253) );
  AOI21_X1 U15375 ( .B1(n13327), .B2(n13270), .A(n13253), .ZN(n13254) );
  OAI21_X1 U15376 ( .B1(n13255), .B2(n15206), .A(n13254), .ZN(P3_U3218) );
  INV_X1 U15377 ( .A(n13256), .ZN(n13259) );
  AOI21_X1 U15378 ( .B1(n13256), .B2(n13257), .A(n13262), .ZN(n13258) );
  AOI21_X1 U15379 ( .B1(n13259), .B2(n14755), .A(n13258), .ZN(n13261) );
  XNOR2_X1 U15380 ( .A(n13261), .B(n13260), .ZN(n13265) );
  AOI22_X1 U15381 ( .A1(n13263), .A2(n15195), .B1(n15192), .B2(n13262), .ZN(
        n13264) );
  OAI21_X1 U15382 ( .B1(n13265), .B2(n15198), .A(n13264), .ZN(n13330) );
  INV_X1 U15383 ( .A(n13330), .ZN(n13272) );
  XNOR2_X1 U15384 ( .A(n6549), .B(n13266), .ZN(n13331) );
  AOI22_X1 U15385 ( .A1(n15206), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15201), 
        .B2(n13267), .ZN(n13268) );
  OAI21_X1 U15386 ( .B1(n15165), .B2(n13385), .A(n13268), .ZN(n13269) );
  AOI21_X1 U15387 ( .B1(n13331), .B2(n13270), .A(n13269), .ZN(n13271) );
  OAI21_X1 U15388 ( .B1(n13272), .B2(n15206), .A(n13271), .ZN(P3_U3219) );
  NOR2_X1 U15389 ( .A1(n15241), .A2(n13335), .ZN(n13274) );
  AOI21_X1 U15390 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n15241), .A(n13274), 
        .ZN(n13273) );
  OAI21_X1 U15391 ( .B1(n13337), .B2(n13334), .A(n13273), .ZN(P3_U3490) );
  AOI21_X1 U15392 ( .B1(P3_REG1_REG_30__SCAN_IN), .B2(n15241), .A(n13274), 
        .ZN(n13275) );
  OAI21_X1 U15393 ( .B1(n13276), .B2(n13334), .A(n13275), .ZN(P3_U3489) );
  NAND2_X1 U15394 ( .A1(n13277), .A2(n13311), .ZN(n13278) );
  OAI211_X1 U15395 ( .C1(n14790), .C2(n13280), .A(n13279), .B(n13278), .ZN(
        n13344) );
  MUX2_X1 U15396 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n13344), .S(n15240), .Z(
        P3_U3487) );
  INV_X1 U15397 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13283) );
  AOI21_X1 U15398 ( .B1(n15223), .B2(n13282), .A(n13281), .ZN(n13345) );
  MUX2_X1 U15399 ( .A(n13283), .B(n13345), .S(n15240), .Z(n13284) );
  OAI21_X1 U15400 ( .B1(n13348), .B2(n13334), .A(n13284), .ZN(P3_U3485) );
  INV_X1 U15401 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13287) );
  AOI21_X1 U15402 ( .B1(n13286), .B2(n14798), .A(n13285), .ZN(n13349) );
  MUX2_X1 U15403 ( .A(n13287), .B(n13349), .S(n15240), .Z(n13288) );
  OAI21_X1 U15404 ( .B1(n13352), .B2(n13334), .A(n13288), .ZN(P3_U3484) );
  INV_X1 U15405 ( .A(n13289), .ZN(n13290) );
  NAND2_X1 U15406 ( .A1(n13290), .A2(n13311), .ZN(n13291) );
  OAI211_X1 U15407 ( .C1(n14790), .C2(n13293), .A(n13292), .B(n13291), .ZN(
        n13353) );
  MUX2_X1 U15408 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13353), .S(n15240), .Z(
        P3_U3483) );
  INV_X1 U15409 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13664) );
  AOI21_X1 U15410 ( .B1(n15223), .B2(n13295), .A(n13294), .ZN(n13354) );
  MUX2_X1 U15411 ( .A(n13664), .B(n13354), .S(n15240), .Z(n13296) );
  OAI21_X1 U15412 ( .B1(n13357), .B2(n13334), .A(n13296), .ZN(P3_U3482) );
  INV_X1 U15413 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13299) );
  AOI21_X1 U15414 ( .B1(n14798), .B2(n13298), .A(n13297), .ZN(n13358) );
  MUX2_X1 U15415 ( .A(n13299), .B(n13358), .S(n15240), .Z(n13300) );
  OAI21_X1 U15416 ( .B1(n13361), .B2(n13334), .A(n13300), .ZN(P3_U3481) );
  INV_X1 U15417 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13303) );
  AOI21_X1 U15418 ( .B1(n13302), .B2(n14798), .A(n13301), .ZN(n13362) );
  MUX2_X1 U15419 ( .A(n13303), .B(n13362), .S(n15240), .Z(n13304) );
  OAI21_X1 U15420 ( .B1(n13365), .B2(n13334), .A(n13304), .ZN(P3_U3480) );
  NAND2_X1 U15421 ( .A1(n13305), .A2(n13311), .ZN(n13306) );
  OAI211_X1 U15422 ( .C1(n14790), .C2(n13308), .A(n13307), .B(n13306), .ZN(
        n13366) );
  MUX2_X1 U15423 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n13366), .S(n15240), .Z(
        P3_U3479) );
  INV_X1 U15424 ( .A(n13309), .ZN(n13312) );
  AOI21_X1 U15425 ( .B1(n13312), .B2(n13311), .A(n13310), .ZN(n13313) );
  OAI21_X1 U15426 ( .B1(n14790), .B2(n13314), .A(n13313), .ZN(n13367) );
  MUX2_X1 U15427 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n13367), .S(n15240), .Z(
        P3_U3478) );
  INV_X1 U15428 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13317) );
  AOI21_X1 U15429 ( .B1(n13316), .B2(n14798), .A(n13315), .ZN(n13368) );
  MUX2_X1 U15430 ( .A(n13317), .B(n13368), .S(n15240), .Z(n13318) );
  OAI21_X1 U15431 ( .B1(n13371), .B2(n13334), .A(n13318), .ZN(P3_U3477) );
  NAND2_X1 U15432 ( .A1(n13319), .A2(n14798), .ZN(n13320) );
  OAI211_X1 U15433 ( .C1(n15226), .C2(n13322), .A(n13321), .B(n13320), .ZN(
        n13372) );
  MUX2_X1 U15434 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13372), .S(n15240), .Z(
        P3_U3476) );
  INV_X1 U15435 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13671) );
  AOI21_X1 U15436 ( .B1(n14798), .B2(n13324), .A(n13323), .ZN(n13373) );
  MUX2_X1 U15437 ( .A(n13671), .B(n13373), .S(n15240), .Z(n13325) );
  OAI21_X1 U15438 ( .B1(n13376), .B2(n13334), .A(n13325), .ZN(P3_U3475) );
  AOI21_X1 U15439 ( .B1(n13327), .B2(n14798), .A(n13326), .ZN(n13377) );
  MUX2_X1 U15440 ( .A(n13328), .B(n13377), .S(n15240), .Z(n13329) );
  OAI21_X1 U15441 ( .B1(n13380), .B2(n13334), .A(n13329), .ZN(P3_U3474) );
  AOI21_X1 U15442 ( .B1(n14798), .B2(n13331), .A(n13330), .ZN(n13381) );
  MUX2_X1 U15443 ( .A(n13332), .B(n13381), .S(n15240), .Z(n13333) );
  OAI21_X1 U15444 ( .B1(n13385), .B2(n13334), .A(n13333), .ZN(P3_U3473) );
  NOR2_X1 U15445 ( .A1(n15234), .A2(n13335), .ZN(n13340) );
  AOI21_X1 U15446 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n15234), .A(n13340), 
        .ZN(n13336) );
  OAI21_X1 U15447 ( .B1(n13337), .B2(n13384), .A(n13336), .ZN(P3_U3458) );
  INV_X1 U15448 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n13343) );
  INV_X1 U15449 ( .A(n13384), .ZN(n13338) );
  NAND2_X1 U15450 ( .A1(n13339), .A2(n13338), .ZN(n13342) );
  INV_X1 U15451 ( .A(n13340), .ZN(n13341) );
  OAI211_X1 U15452 ( .C1(n13343), .C2(n15232), .A(n13342), .B(n13341), .ZN(
        P3_U3457) );
  MUX2_X1 U15453 ( .A(P3_REG0_REG_28__SCAN_IN), .B(n13344), .S(n15232), .Z(
        P3_U3455) );
  INV_X1 U15454 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13346) );
  MUX2_X1 U15455 ( .A(n13346), .B(n13345), .S(n15232), .Z(n13347) );
  OAI21_X1 U15456 ( .B1(n13348), .B2(n13384), .A(n13347), .ZN(P3_U3453) );
  INV_X1 U15457 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13350) );
  MUX2_X1 U15458 ( .A(n13350), .B(n13349), .S(n15232), .Z(n13351) );
  OAI21_X1 U15459 ( .B1(n13352), .B2(n13384), .A(n13351), .ZN(P3_U3452) );
  MUX2_X1 U15460 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n13353), .S(n15232), .Z(
        P3_U3451) );
  INV_X1 U15461 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13355) );
  MUX2_X1 U15462 ( .A(n13355), .B(n13354), .S(n15232), .Z(n13356) );
  OAI21_X1 U15463 ( .B1(n13357), .B2(n13384), .A(n13356), .ZN(P3_U3450) );
  INV_X1 U15464 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13359) );
  MUX2_X1 U15465 ( .A(n13359), .B(n13358), .S(n15232), .Z(n13360) );
  OAI21_X1 U15466 ( .B1(n13361), .B2(n13384), .A(n13360), .ZN(P3_U3449) );
  INV_X1 U15467 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13363) );
  MUX2_X1 U15468 ( .A(n13363), .B(n13362), .S(n15232), .Z(n13364) );
  OAI21_X1 U15469 ( .B1(n13365), .B2(n13384), .A(n13364), .ZN(P3_U3448) );
  MUX2_X1 U15470 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n13366), .S(n15232), .Z(
        P3_U3447) );
  MUX2_X1 U15471 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n13367), .S(n15232), .Z(
        P3_U3446) );
  INV_X1 U15472 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13369) );
  MUX2_X1 U15473 ( .A(n13369), .B(n13368), .S(n15232), .Z(n13370) );
  OAI21_X1 U15474 ( .B1(n13371), .B2(n13384), .A(n13370), .ZN(P3_U3444) );
  MUX2_X1 U15475 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n13372), .S(n15232), .Z(
        P3_U3441) );
  INV_X1 U15476 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13374) );
  MUX2_X1 U15477 ( .A(n13374), .B(n13373), .S(n15232), .Z(n13375) );
  OAI21_X1 U15478 ( .B1(n13376), .B2(n13384), .A(n13375), .ZN(P3_U3438) );
  INV_X1 U15479 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13378) );
  MUX2_X1 U15480 ( .A(n13378), .B(n13377), .S(n15232), .Z(n13379) );
  OAI21_X1 U15481 ( .B1(n13380), .B2(n13384), .A(n13379), .ZN(P3_U3435) );
  INV_X1 U15482 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13382) );
  MUX2_X1 U15483 ( .A(n13382), .B(n13381), .S(n15232), .Z(n13383) );
  OAI21_X1 U15484 ( .B1(n13385), .B2(n13384), .A(n13383), .ZN(P3_U3432) );
  MUX2_X1 U15485 ( .A(P3_D_REG_1__SCAN_IN), .B(n13386), .S(n13387), .Z(
        P3_U3377) );
  MUX2_X1 U15486 ( .A(P3_D_REG_0__SCAN_IN), .B(n13388), .S(n13387), .Z(
        P3_U3376) );
  INV_X1 U15487 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13389) );
  NAND3_X1 U15488 ( .A1(n13389), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n13391) );
  OAI22_X1 U15489 ( .A1(n7612), .A2(n13391), .B1(n13390), .B2(n9579), .ZN(
        n13392) );
  AOI21_X1 U15490 ( .B1(n13394), .B2(n13393), .A(n13392), .ZN(n13395) );
  INV_X1 U15491 ( .A(n13395), .ZN(P3_U3264) );
  INV_X1 U15492 ( .A(n13396), .ZN(n13398) );
  OAI222_X1 U15493 ( .A1(n9579), .A2(n13399), .B1(n12508), .B2(n13398), .C1(
        n13397), .C2(P3_U3151), .ZN(P3_U3266) );
  INV_X1 U15494 ( .A(n13400), .ZN(n13401) );
  OAI222_X1 U15495 ( .A1(n9579), .A2(n13402), .B1(P3_U3151), .B2(n8044), .C1(
        n12508), .C2(n13401), .ZN(P3_U3267) );
  NOR3_X1 U15496 ( .A1(n13512), .A2(n13404), .A3(n13403), .ZN(n13410) );
  AOI21_X1 U15497 ( .B1(n13406), .B2(n13405), .A(n13478), .ZN(n13409) );
  INV_X1 U15498 ( .A(n13407), .ZN(n13408) );
  OAI21_X1 U15499 ( .B1(n13410), .B2(n13409), .A(n13408), .ZN(n13418) );
  INV_X1 U15500 ( .A(n13411), .ZN(n13412) );
  OAI22_X1 U15501 ( .A1(n13503), .A2(n13412), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13710), .ZN(n13413) );
  INV_X1 U15502 ( .A(n13413), .ZN(n13417) );
  NAND2_X1 U15503 ( .A1(n13522), .A2(n15063), .ZN(n13416) );
  NAND2_X1 U15504 ( .A1(n13510), .A2(n13414), .ZN(n13415) );
  NAND4_X1 U15505 ( .A1(n13418), .A2(n13417), .A3(n13416), .A4(n13415), .ZN(
        P2_U3185) );
  INV_X1 U15506 ( .A(n13954), .ZN(n13434) );
  INV_X1 U15507 ( .A(n13419), .ZN(n13420) );
  XNOR2_X1 U15508 ( .A(n13960), .B(n13424), .ZN(n13423) );
  NAND2_X1 U15509 ( .A1(n13536), .A2(n6649), .ZN(n13422) );
  XNOR2_X1 U15510 ( .A(n13423), .B(n13422), .ZN(n13516) );
  XNOR2_X1 U15511 ( .A(n13954), .B(n13424), .ZN(n13426) );
  NAND2_X1 U15512 ( .A1(n13535), .A2(n13845), .ZN(n13425) );
  NOR2_X1 U15513 ( .A1(n13426), .A2(n13425), .ZN(n13456) );
  AOI21_X1 U15514 ( .B1(n13426), .B2(n13425), .A(n13456), .ZN(n13427) );
  OAI211_X1 U15515 ( .C1(n6503), .C2(n13427), .A(n13458), .B(n13527), .ZN(
        n13433) );
  NAND2_X1 U15516 ( .A1(n13534), .A2(n13517), .ZN(n13429) );
  NAND2_X1 U15517 ( .A1(n13536), .A2(n13518), .ZN(n13428) );
  NAND2_X1 U15518 ( .A1(n13429), .A2(n13428), .ZN(n13760) );
  OAI22_X1 U15519 ( .A1(n13763), .A2(n13495), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13430), .ZN(n13431) );
  AOI21_X1 U15520 ( .B1(n13760), .B2(n13521), .A(n13431), .ZN(n13432) );
  OAI211_X1 U15521 ( .C1(n13434), .C2(n13525), .A(n13433), .B(n13432), .ZN(
        P2_U3186) );
  INV_X1 U15522 ( .A(n13435), .ZN(n13443) );
  AOI22_X1 U15523 ( .A1(n13437), .A2(n13527), .B1(n13436), .B2(n13539), .ZN(
        n13442) );
  AOI22_X1 U15524 ( .A1(n13538), .A2(n13517), .B1(n13518), .B2(n13540), .ZN(
        n13821) );
  INV_X1 U15525 ( .A(n13821), .ZN(n13438) );
  AOI22_X1 U15526 ( .A1(n13438), .A2(n13521), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13439) );
  OAI21_X1 U15527 ( .B1(n13824), .B2(n13495), .A(n13439), .ZN(n13440) );
  AOI21_X1 U15528 ( .B1(n13977), .B2(n13510), .A(n13440), .ZN(n13441) );
  OAI21_X1 U15529 ( .B1(n13443), .B2(n13442), .A(n13441), .ZN(P2_U3188) );
  INV_X1 U15530 ( .A(n13444), .ZN(n13505) );
  NOR3_X1 U15531 ( .A1(n13446), .A2(n13445), .A3(n13512), .ZN(n13447) );
  AOI21_X1 U15532 ( .B1(n13505), .B2(n13527), .A(n13447), .ZN(n13455) );
  INV_X1 U15533 ( .A(n6424), .ZN(n13452) );
  AND2_X1 U15534 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13577) );
  AOI22_X1 U15535 ( .A1(n13542), .A2(n13517), .B1(n13518), .B2(n13544), .ZN(
        n13893) );
  NOR2_X1 U15536 ( .A1(n13503), .A2(n13893), .ZN(n13449) );
  AOI211_X1 U15537 ( .C1(n13522), .C2(n13900), .A(n13577), .B(n13449), .ZN(
        n13450) );
  OAI21_X1 U15538 ( .B1(n14059), .B2(n13525), .A(n13450), .ZN(n13451) );
  AOI21_X1 U15539 ( .B1(n13452), .B2(n13527), .A(n13451), .ZN(n13453) );
  OAI21_X1 U15540 ( .B1(n13455), .B2(n13454), .A(n13453), .ZN(P2_U3191) );
  INV_X1 U15541 ( .A(n13456), .ZN(n13457) );
  NAND2_X1 U15542 ( .A1(n13458), .A2(n13457), .ZN(n13463) );
  NAND2_X1 U15543 ( .A1(n13534), .A2(n13845), .ZN(n13460) );
  XNOR2_X1 U15544 ( .A(n13460), .B(n6627), .ZN(n13461) );
  XNOR2_X1 U15545 ( .A(n13608), .B(n13461), .ZN(n13462) );
  XNOR2_X1 U15546 ( .A(n13463), .B(n13462), .ZN(n13470) );
  NOR2_X1 U15547 ( .A1(n13602), .A2(n13495), .ZN(n13468) );
  NAND2_X1 U15548 ( .A1(n13533), .A2(n13517), .ZN(n13465) );
  NAND2_X1 U15549 ( .A1(n13535), .A2(n13518), .ZN(n13464) );
  AND2_X1 U15550 ( .A1(n13465), .A2(n13464), .ZN(n13594) );
  OAI22_X1 U15551 ( .A1(n13594), .A2(n13503), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13466), .ZN(n13467) );
  AOI211_X1 U15552 ( .C1(n13608), .C2(n13510), .A(n13468), .B(n13467), .ZN(
        n13469) );
  OAI21_X1 U15553 ( .B1(n13470), .B2(n13478), .A(n13469), .ZN(P2_U3192) );
  XNOR2_X1 U15554 ( .A(n6764), .B(n13471), .ZN(n13472) );
  XNOR2_X1 U15555 ( .A(n13473), .B(n13472), .ZN(n13479) );
  AOI22_X1 U15556 ( .A1(n13540), .A2(n13517), .B1(n13518), .B2(n13542), .ZN(
        n13859) );
  OAI22_X1 U15557 ( .A1(n13859), .A2(n13503), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13474), .ZN(n13475) );
  AOI21_X1 U15558 ( .B1(n13863), .B2(n13522), .A(n13475), .ZN(n13477) );
  NAND2_X1 U15559 ( .A1(n14050), .A2(n13510), .ZN(n13476) );
  OAI211_X1 U15560 ( .C1(n13479), .C2(n13478), .A(n13477), .B(n13476), .ZN(
        P2_U3195) );
  OAI211_X1 U15561 ( .C1(n13482), .C2(n13481), .A(n13480), .B(n13527), .ZN(
        n13488) );
  NAND2_X1 U15562 ( .A1(n13537), .A2(n13517), .ZN(n13484) );
  NAND2_X1 U15563 ( .A1(n13539), .A2(n13518), .ZN(n13483) );
  NAND2_X1 U15564 ( .A1(n13484), .A2(n13483), .ZN(n13807) );
  AOI22_X1 U15565 ( .A1(n13807), .A2(n13521), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13485) );
  OAI21_X1 U15566 ( .B1(n13811), .B2(n13495), .A(n13485), .ZN(n13486) );
  AOI21_X1 U15567 ( .B1(n13973), .B2(n13510), .A(n13486), .ZN(n13487) );
  NAND2_X1 U15568 ( .A1(n13488), .A2(n13487), .ZN(P2_U3201) );
  NAND2_X1 U15569 ( .A1(n13490), .A2(n13489), .ZN(n13492) );
  XOR2_X1 U15570 ( .A(n13492), .B(n13491), .Z(n13498) );
  AOI22_X1 U15571 ( .A1(n13541), .A2(n13517), .B1(n13518), .B2(n13543), .ZN(
        n13874) );
  INV_X1 U15572 ( .A(n13874), .ZN(n13493) );
  AOI22_X1 U15573 ( .A1(n13493), .A2(n13521), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13494) );
  OAI21_X1 U15574 ( .B1(n13882), .B2(n13495), .A(n13494), .ZN(n13496) );
  AOI21_X1 U15575 ( .B1(n13881), .B2(n13510), .A(n13496), .ZN(n13497) );
  OAI21_X1 U15576 ( .B1(n13498), .B2(n13478), .A(n13497), .ZN(P2_U3205) );
  INV_X1 U15577 ( .A(n13499), .ZN(n13500) );
  NAND2_X1 U15578 ( .A1(n13522), .A2(n13500), .ZN(n13502) );
  OAI211_X1 U15579 ( .C1(n13504), .C2(n13503), .A(n13502), .B(n13501), .ZN(
        n13509) );
  AOI211_X1 U15580 ( .C1(n13507), .C2(n13506), .A(n13478), .B(n13505), .ZN(
        n13508) );
  AOI211_X1 U15581 ( .C1(n14006), .C2(n13510), .A(n13509), .B(n13508), .ZN(
        n13511) );
  INV_X1 U15582 ( .A(n13511), .ZN(P2_U3210) );
  NOR3_X1 U15583 ( .A1(n13514), .A2(n13513), .A3(n13512), .ZN(n13515) );
  AOI21_X1 U15584 ( .B1(n13421), .B2(n13527), .A(n13515), .ZN(n13531) );
  INV_X1 U15585 ( .A(n13516), .ZN(n13530) );
  NAND2_X1 U15586 ( .A1(n13535), .A2(n13517), .ZN(n13520) );
  NAND2_X1 U15587 ( .A1(n13537), .A2(n13518), .ZN(n13519) );
  NAND2_X1 U15588 ( .A1(n13520), .A2(n13519), .ZN(n13773) );
  AOI22_X1 U15589 ( .A1(n13773), .A2(n13521), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13524) );
  NAND2_X1 U15590 ( .A1(n13778), .A2(n13522), .ZN(n13523) );
  OAI211_X1 U15591 ( .C1(n13780), .C2(n13525), .A(n13524), .B(n13523), .ZN(
        n13526) );
  AOI21_X1 U15592 ( .B1(n13528), .B2(n13527), .A(n13526), .ZN(n13529) );
  OAI21_X1 U15593 ( .B1(n13531), .B2(n13530), .A(n13529), .ZN(P2_U3212) );
  MUX2_X1 U15594 ( .A(n13581), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13562), .Z(
        P2_U3562) );
  MUX2_X1 U15595 ( .A(n13532), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13562), .Z(
        P2_U3561) );
  MUX2_X1 U15596 ( .A(n13533), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13562), .Z(
        P2_U3560) );
  MUX2_X1 U15597 ( .A(n13534), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13562), .Z(
        P2_U3559) );
  MUX2_X1 U15598 ( .A(n13535), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13562), .Z(
        P2_U3558) );
  MUX2_X1 U15599 ( .A(n13536), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13562), .Z(
        P2_U3557) );
  MUX2_X1 U15600 ( .A(n13537), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13562), .Z(
        P2_U3556) );
  MUX2_X1 U15601 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13538), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15602 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13539), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U15603 ( .A(n13540), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13562), .Z(
        P2_U3553) );
  MUX2_X1 U15604 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13541), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15605 ( .A(n13542), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13562), .Z(
        P2_U3551) );
  MUX2_X1 U15606 ( .A(n13543), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13562), .Z(
        P2_U3550) );
  MUX2_X1 U15607 ( .A(n13544), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13562), .Z(
        P2_U3549) );
  MUX2_X1 U15608 ( .A(n13545), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13562), .Z(
        P2_U3548) );
  MUX2_X1 U15609 ( .A(n13546), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13562), .Z(
        P2_U3547) );
  MUX2_X1 U15610 ( .A(n13547), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13562), .Z(
        P2_U3546) );
  MUX2_X1 U15611 ( .A(n13548), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13562), .Z(
        P2_U3545) );
  MUX2_X1 U15612 ( .A(n13549), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13562), .Z(
        P2_U3544) );
  MUX2_X1 U15613 ( .A(n13550), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13562), .Z(
        P2_U3543) );
  MUX2_X1 U15614 ( .A(n13551), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13562), .Z(
        P2_U3542) );
  MUX2_X1 U15615 ( .A(n13552), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13562), .Z(
        P2_U3541) );
  MUX2_X1 U15616 ( .A(n13553), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13562), .Z(
        P2_U3540) );
  MUX2_X1 U15617 ( .A(n13554), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13562), .Z(
        P2_U3539) );
  MUX2_X1 U15618 ( .A(n13555), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13562), .Z(
        P2_U3538) );
  MUX2_X1 U15619 ( .A(n13556), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13562), .Z(
        P2_U3537) );
  MUX2_X1 U15620 ( .A(n13557), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13562), .Z(
        P2_U3536) );
  MUX2_X1 U15621 ( .A(n13558), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13562), .Z(
        P2_U3535) );
  MUX2_X1 U15622 ( .A(n13559), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13562), .Z(
        P2_U3534) );
  MUX2_X1 U15623 ( .A(n13560), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13562), .Z(
        P2_U3533) );
  MUX2_X1 U15624 ( .A(n13561), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13562), .Z(
        P2_U3532) );
  MUX2_X1 U15625 ( .A(n13563), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13562), .Z(
        P2_U3531) );
  NOR2_X1 U15626 ( .A1(n13565), .A2(n13564), .ZN(n13566) );
  XNOR2_X1 U15627 ( .A(n13566), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13571) );
  NOR2_X1 U15628 ( .A1(n13568), .A2(n13567), .ZN(n13569) );
  INV_X1 U15629 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13684) );
  XOR2_X1 U15630 ( .A(n13569), .B(n13684), .Z(n13573) );
  NAND2_X1 U15631 ( .A1(n13573), .A2(n15039), .ZN(n13570) );
  INV_X1 U15632 ( .A(n13571), .ZN(n13572) );
  OAI22_X1 U15633 ( .A1(n13573), .A2(n15054), .B1(n13572), .B2(n15046), .ZN(
        n13575) );
  INV_X1 U15634 ( .A(n13578), .ZN(P2_U3233) );
  NAND2_X1 U15635 ( .A1(n14028), .A2(n13586), .ZN(n13585) );
  XNOR2_X1 U15636 ( .A(n13579), .B(n13585), .ZN(n13580) );
  NAND2_X1 U15637 ( .A1(n13934), .A2(n15064), .ZN(n13584) );
  AND2_X1 U15638 ( .A1(n13582), .A2(n13581), .ZN(n13933) );
  INV_X1 U15639 ( .A(n13933), .ZN(n13937) );
  NOR2_X1 U15640 ( .A1(n15075), .A2(n13937), .ZN(n13588) );
  AOI21_X1 U15641 ( .B1(n15075), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13588), 
        .ZN(n13583) );
  OAI211_X1 U15642 ( .C1(n14024), .C2(n15069), .A(n13584), .B(n13583), .ZN(
        P2_U3234) );
  OAI211_X1 U15643 ( .C1(n14028), .C2(n13586), .A(n9326), .B(n13585), .ZN(
        n13938) );
  NOR2_X1 U15644 ( .A1(n14028), .A2(n15069), .ZN(n13587) );
  AOI211_X1 U15645 ( .C1(n15075), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13588), 
        .B(n13587), .ZN(n13589) );
  OAI21_X1 U15646 ( .B1(n13866), .B2(n13938), .A(n13589), .ZN(P2_U3235) );
  NAND3_X1 U15647 ( .A1(n13593), .A2(n13891), .A3(n13592), .ZN(n13595) );
  NAND2_X1 U15648 ( .A1(n13595), .A2(n13594), .ZN(n13948) );
  AOI21_X1 U15649 ( .B1(n13608), .B2(n13765), .A(n6649), .ZN(n13600) );
  OAI22_X1 U15650 ( .A1(n6485), .A2(n13603), .B1(n13825), .B2(n13602), .ZN(
        n13604) );
  OAI21_X1 U15651 ( .B1(n13948), .B2(n13607), .A(n13868), .ZN(n13611) );
  NAND2_X1 U15652 ( .A1(n13949), .A2(n13925), .ZN(n13610) );
  AOI22_X1 U15653 ( .A1(n13608), .A2(n13927), .B1(n15075), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n13609) );
  NAND2_X1 U15654 ( .A1(n13611), .A2(n7419), .ZN(n13757) );
  INV_X1 U15655 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n14915) );
  AOI22_X1 U15656 ( .A1(n14915), .A2(keyinput4), .B1(keyinput9), .B2(n13613), 
        .ZN(n13612) );
  OAI221_X1 U15657 ( .B1(n14915), .B2(keyinput4), .C1(n13613), .C2(keyinput9), 
        .A(n13612), .ZN(n13626) );
  AOI22_X1 U15658 ( .A1(n13616), .A2(keyinput34), .B1(n13615), .B2(keyinput50), 
        .ZN(n13614) );
  OAI221_X1 U15659 ( .B1(n13616), .B2(keyinput34), .C1(n13615), .C2(keyinput50), .A(n13614), .ZN(n13625) );
  AOI22_X1 U15660 ( .A1(n13619), .A2(keyinput22), .B1(n13618), .B2(keyinput63), 
        .ZN(n13617) );
  OAI221_X1 U15661 ( .B1(n13619), .B2(keyinput22), .C1(n13618), .C2(keyinput63), .A(n13617), .ZN(n13624) );
  INV_X1 U15662 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n13621) );
  AOI22_X1 U15663 ( .A1(n13622), .A2(keyinput5), .B1(n13621), .B2(keyinput58), 
        .ZN(n13620) );
  OAI221_X1 U15664 ( .B1(n13622), .B2(keyinput5), .C1(n13621), .C2(keyinput58), 
        .A(n13620), .ZN(n13623) );
  OR4_X1 U15665 ( .A1(n13626), .A2(n13625), .A3(n13624), .A4(n13623), .ZN(
        n13681) );
  AOI22_X1 U15666 ( .A1(n13762), .A2(keyinput0), .B1(n13726), .B2(keyinput7), 
        .ZN(n13627) );
  OAI221_X1 U15667 ( .B1(n13762), .B2(keyinput0), .C1(n13726), .C2(keyinput7), 
        .A(n13627), .ZN(n13630) );
  INV_X1 U15668 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n15078) );
  AOI22_X1 U15669 ( .A1(n15078), .A2(keyinput32), .B1(keyinput37), .B2(n14596), 
        .ZN(n13628) );
  OAI221_X1 U15670 ( .B1(n15078), .B2(keyinput32), .C1(n14596), .C2(keyinput37), .A(n13628), .ZN(n13629) );
  NOR2_X1 U15671 ( .A1(n13630), .A2(n13629), .ZN(n13651) );
  AOI22_X1 U15672 ( .A1(n13632), .A2(keyinput35), .B1(keyinput55), .B2(n13742), 
        .ZN(n13631) );
  OAI221_X1 U15673 ( .B1(n13632), .B2(keyinput35), .C1(n13742), .C2(keyinput55), .A(n13631), .ZN(n13636) );
  INV_X1 U15674 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14187) );
  AOI22_X1 U15675 ( .A1(n14187), .A2(keyinput53), .B1(keyinput61), .B2(n13634), 
        .ZN(n13633) );
  OAI221_X1 U15676 ( .B1(n14187), .B2(keyinput53), .C1(n13634), .C2(keyinput61), .A(n13633), .ZN(n13635) );
  NOR2_X1 U15677 ( .A1(n13636), .A2(n13635), .ZN(n13650) );
  INV_X1 U15678 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n14913) );
  INV_X1 U15679 ( .A(keyinput20), .ZN(n13637) );
  XNOR2_X1 U15680 ( .A(n14913), .B(n13637), .ZN(n13649) );
  XNOR2_X1 U15681 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(keyinput30), .ZN(n13641)
         );
  XNOR2_X1 U15682 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput24), .ZN(n13640) );
  XNOR2_X1 U15683 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput33), .ZN(n13639) );
  XNOR2_X1 U15684 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput13), .ZN(n13638) );
  NAND4_X1 U15685 ( .A1(n13641), .A2(n13640), .A3(n13639), .A4(n13638), .ZN(
        n13647) );
  XNOR2_X1 U15686 ( .A(P2_REG1_REG_13__SCAN_IN), .B(keyinput1), .ZN(n13645) );
  XNOR2_X1 U15687 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput3), .ZN(n13644) );
  XNOR2_X1 U15688 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput51), .ZN(n13643) );
  XNOR2_X1 U15689 ( .A(keyinput19), .B(P2_REG3_REG_13__SCAN_IN), .ZN(n13642)
         );
  NAND4_X1 U15690 ( .A1(n13645), .A2(n13644), .A3(n13643), .A4(n13642), .ZN(
        n13646) );
  NOR2_X1 U15691 ( .A1(n13647), .A2(n13646), .ZN(n13648) );
  NAND4_X1 U15692 ( .A1(n13651), .A2(n13650), .A3(n13649), .A4(n13648), .ZN(
        n13680) );
  AOI22_X1 U15693 ( .A1(n13653), .A2(keyinput17), .B1(n13735), .B2(keyinput27), 
        .ZN(n13652) );
  OAI221_X1 U15694 ( .B1(n13653), .B2(keyinput17), .C1(n13735), .C2(keyinput27), .A(n13652), .ZN(n13658) );
  AOI22_X1 U15695 ( .A1(n9157), .A2(keyinput38), .B1(n13655), .B2(keyinput42), 
        .ZN(n13654) );
  OAI221_X1 U15696 ( .B1(n9157), .B2(keyinput38), .C1(n13655), .C2(keyinput42), 
        .A(n13654), .ZN(n13657) );
  INV_X1 U15697 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15077) );
  XNOR2_X1 U15698 ( .A(n15077), .B(keyinput41), .ZN(n13656) );
  NOR3_X1 U15699 ( .A1(n13658), .A2(n13657), .A3(n13656), .ZN(n13678) );
  AOI22_X1 U15700 ( .A1(n13661), .A2(keyinput16), .B1(keyinput8), .B2(n13660), 
        .ZN(n13659) );
  OAI221_X1 U15701 ( .B1(n13661), .B2(keyinput16), .C1(n13660), .C2(keyinput8), 
        .A(n13659), .ZN(n13669) );
  INV_X1 U15702 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n13663) );
  AOI22_X1 U15703 ( .A1(n13664), .A2(keyinput56), .B1(n13663), .B2(keyinput54), 
        .ZN(n13662) );
  OAI221_X1 U15704 ( .B1(n13664), .B2(keyinput56), .C1(n13663), .C2(keyinput54), .A(n13662), .ZN(n13668) );
  INV_X1 U15705 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n13666) );
  AOI22_X1 U15706 ( .A1(n13666), .A2(keyinput25), .B1(n14087), .B2(keyinput11), 
        .ZN(n13665) );
  OAI221_X1 U15707 ( .B1(n13666), .B2(keyinput25), .C1(n14087), .C2(keyinput11), .A(n13665), .ZN(n13667) );
  NOR3_X1 U15708 ( .A1(n13669), .A2(n13668), .A3(n13667), .ZN(n13677) );
  AOI22_X1 U15709 ( .A1(n13671), .A2(keyinput59), .B1(keyinput26), .B2(n8787), 
        .ZN(n13670) );
  OAI221_X1 U15710 ( .B1(n13671), .B2(keyinput59), .C1(n8787), .C2(keyinput26), 
        .A(n13670), .ZN(n13675) );
  AOI22_X1 U15711 ( .A1(n8495), .A2(keyinput48), .B1(keyinput21), .B2(n13673), 
        .ZN(n13672) );
  OAI221_X1 U15712 ( .B1(n8495), .B2(keyinput48), .C1(n13673), .C2(keyinput21), 
        .A(n13672), .ZN(n13674) );
  NOR2_X1 U15713 ( .A1(n13675), .A2(n13674), .ZN(n13676) );
  NAND3_X1 U15714 ( .A1(n13678), .A2(n13677), .A3(n13676), .ZN(n13679) );
  NOR3_X1 U15715 ( .A1(n13681), .A2(n13680), .A3(n13679), .ZN(n13722) );
  AOI22_X1 U15716 ( .A1(n13684), .A2(keyinput12), .B1(keyinput29), .B2(n13683), 
        .ZN(n13682) );
  OAI221_X1 U15717 ( .B1(n13684), .B2(keyinput12), .C1(n13683), .C2(keyinput29), .A(n13682), .ZN(n13695) );
  AOI22_X1 U15718 ( .A1(n13687), .A2(keyinput23), .B1(keyinput18), .B2(n13686), 
        .ZN(n13685) );
  OAI221_X1 U15719 ( .B1(n13687), .B2(keyinput23), .C1(n13686), .C2(keyinput18), .A(n13685), .ZN(n13694) );
  AOI22_X1 U15720 ( .A1(n13741), .A2(keyinput57), .B1(n13689), .B2(keyinput47), 
        .ZN(n13688) );
  OAI221_X1 U15721 ( .B1(n13741), .B2(keyinput57), .C1(n13689), .C2(keyinput47), .A(n13688), .ZN(n13693) );
  INV_X1 U15722 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n14914) );
  INV_X1 U15723 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13691) );
  AOI22_X1 U15724 ( .A1(n14914), .A2(keyinput43), .B1(n13691), .B2(keyinput46), 
        .ZN(n13690) );
  OAI221_X1 U15725 ( .B1(n14914), .B2(keyinput43), .C1(n13691), .C2(keyinput46), .A(n13690), .ZN(n13692) );
  NOR4_X1 U15726 ( .A1(n13695), .A2(n13694), .A3(n13693), .A4(n13692), .ZN(
        n13721) );
  INV_X1 U15727 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n13697) );
  AOI22_X1 U15728 ( .A1(n13740), .A2(keyinput31), .B1(keyinput10), .B2(n13697), 
        .ZN(n13696) );
  OAI221_X1 U15729 ( .B1(n13740), .B2(keyinput31), .C1(n13697), .C2(keyinput10), .A(n13696), .ZN(n13707) );
  INV_X1 U15730 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n13699) );
  AOI22_X1 U15731 ( .A1(n13727), .A2(keyinput14), .B1(keyinput44), .B2(n13699), 
        .ZN(n13698) );
  OAI221_X1 U15732 ( .B1(n13727), .B2(keyinput14), .C1(n13699), .C2(keyinput44), .A(n13698), .ZN(n13706) );
  INV_X1 U15733 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n15079) );
  AOI22_X1 U15734 ( .A1(n13701), .A2(keyinput28), .B1(n15079), .B2(keyinput39), 
        .ZN(n13700) );
  OAI221_X1 U15735 ( .B1(n13701), .B2(keyinput28), .C1(n15079), .C2(keyinput39), .A(n13700), .ZN(n13705) );
  INV_X1 U15736 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n13703) );
  AOI22_X1 U15737 ( .A1(n13703), .A2(keyinput60), .B1(keyinput52), .B2(n14112), 
        .ZN(n13702) );
  OAI221_X1 U15738 ( .B1(n13703), .B2(keyinput60), .C1(n14112), .C2(keyinput52), .A(n13702), .ZN(n13704) );
  NOR4_X1 U15739 ( .A1(n13707), .A2(n13706), .A3(n13705), .A4(n13704), .ZN(
        n13720) );
  AOI22_X1 U15740 ( .A1(n13710), .A2(keyinput45), .B1(keyinput40), .B2(n13709), 
        .ZN(n13708) );
  OAI221_X1 U15741 ( .B1(n13710), .B2(keyinput45), .C1(n13709), .C2(keyinput40), .A(n13708), .ZN(n13718) );
  AOI22_X1 U15742 ( .A1(n10945), .A2(keyinput6), .B1(n13731), .B2(keyinput36), 
        .ZN(n13711) );
  OAI221_X1 U15743 ( .B1(n10945), .B2(keyinput6), .C1(n13731), .C2(keyinput36), 
        .A(n13711), .ZN(n13717) );
  AOI22_X1 U15744 ( .A1(n13725), .A2(keyinput49), .B1(keyinput2), .B2(n6807), 
        .ZN(n13712) );
  OAI221_X1 U15745 ( .B1(n13725), .B2(keyinput49), .C1(n6807), .C2(keyinput2), 
        .A(n13712), .ZN(n13716) );
  AOI22_X1 U15746 ( .A1(n13714), .A2(keyinput62), .B1(n14484), .B2(keyinput15), 
        .ZN(n13713) );
  OAI221_X1 U15747 ( .B1(n13714), .B2(keyinput62), .C1(n14484), .C2(keyinput15), .A(n13713), .ZN(n13715) );
  NOR4_X1 U15748 ( .A1(n13718), .A2(n13717), .A3(n13716), .A4(n13715), .ZN(
        n13719) );
  NAND4_X1 U15749 ( .A1(n13722), .A2(n13721), .A3(n13720), .A4(n13719), .ZN(
        n13755) );
  NOR4_X1 U15750 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_REG1_REG_4__SCAN_IN), 
        .A3(P1_ADDR_REG_14__SCAN_IN), .A4(P3_DATAO_REG_29__SCAN_IN), .ZN(
        n13723) );
  NAND4_X1 U15751 ( .A1(n13724), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_REG0_REG_2__SCAN_IN), .A4(n13723), .ZN(n13739) );
  NAND4_X1 U15752 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), 
        .A3(P2_REG3_REG_12__SCAN_IN), .A4(n13762), .ZN(n13738) );
  NAND4_X1 U15753 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(P2_REG2_REG_16__SCAN_IN), 
        .A3(P2_REG2_REG_11__SCAN_IN), .A4(n13725), .ZN(n13730) );
  NAND4_X1 U15754 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(SI_16_), .A3(n14087), 
        .A4(n13726), .ZN(n13729) );
  NAND4_X1 U15755 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .A3(n10426), .A4(n13727), .ZN(n13728) );
  NOR4_X1 U15756 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n13730), .A3(n13729), 
        .A4(n13728), .ZN(n13733) );
  NAND4_X1 U15757 ( .A1(n13733), .A2(P2_REG2_REG_19__SCAN_IN), .A3(n13732), 
        .A4(n13731), .ZN(n13737) );
  NAND4_X1 U15758 ( .A1(n13735), .A2(n13734), .A3(P2_DATAO_REG_21__SCAN_IN), 
        .A4(P2_IR_REG_26__SCAN_IN), .ZN(n13736) );
  NOR4_X1 U15759 ( .A1(n13739), .A2(n13738), .A3(n13737), .A4(n13736), .ZN(
        n13753) );
  NAND4_X1 U15760 ( .A1(n13741), .A2(n13740), .A3(n14913), .A4(n8787), .ZN(
        n13745) );
  NAND3_X1 U15761 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_REG3_REG_24__SCAN_IN), 
        .A3(n13742), .ZN(n13744) );
  NAND4_X1 U15762 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .A3(P3_ADDR_REG_15__SCAN_IN), .A4(P3_DATAO_REG_27__SCAN_IN), .ZN(
        n13743) );
  NOR4_X1 U15763 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(n13745), .A3(n13744), 
        .A4(n13743), .ZN(n13752) );
  NAND4_X1 U15764 ( .A1(P3_D_REG_10__SCAN_IN), .A2(P3_D_REG_7__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_DATAO_REG_3__SCAN_IN), .ZN(n13749) );
  NAND4_X1 U15765 ( .A1(P1_REG0_REG_27__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .A3(P1_REG3_REG_14__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n13748)
         );
  NAND4_X1 U15766 ( .A1(P3_REG1_REG_24__SCAN_IN), .A2(P3_REG1_REG_23__SCAN_IN), 
        .A3(P1_REG2_REG_31__SCAN_IN), .A4(P2_ADDR_REG_11__SCAN_IN), .ZN(n13747) );
  NAND4_X1 U15767 ( .A1(P3_REG2_REG_28__SCAN_IN), .A2(P3_REG2_REG_18__SCAN_IN), 
        .A3(P3_REG1_REG_16__SCAN_IN), .A4(P3_REG2_REG_31__SCAN_IN), .ZN(n13746) );
  NOR4_X1 U15768 ( .A1(n13749), .A2(n13748), .A3(n13747), .A4(n13746), .ZN(
        n13751) );
  NOR4_X1 U15769 ( .A1(P1_REG1_REG_24__SCAN_IN), .A2(P1_REG2_REG_19__SCAN_IN), 
        .A3(P1_REG0_REG_18__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n13750) );
  NAND4_X1 U15770 ( .A1(n13753), .A2(n13752), .A3(n13751), .A4(n13750), .ZN(
        n13754) );
  XNOR2_X1 U15771 ( .A(n13755), .B(n13754), .ZN(n13756) );
  XNOR2_X1 U15772 ( .A(n13757), .B(n13756), .ZN(P2_U3237) );
  XNOR2_X1 U15773 ( .A(n13759), .B(n13758), .ZN(n13761) );
  AOI21_X1 U15774 ( .B1(n13761), .B2(n13891), .A(n13760), .ZN(n13957) );
  OAI22_X1 U15775 ( .A1(n13763), .A2(n13825), .B1(n13762), .B2(n13868), .ZN(
        n13767) );
  NAND2_X1 U15776 ( .A1(n13954), .A2(n13775), .ZN(n13764) );
  NAND3_X1 U15777 ( .A1(n13765), .A2(n9326), .A3(n13764), .ZN(n13955) );
  NOR2_X1 U15778 ( .A1(n13955), .A2(n13866), .ZN(n13766) );
  AOI211_X1 U15779 ( .C1(n13927), .C2(n13954), .A(n13767), .B(n13766), .ZN(
        n13771) );
  OR2_X1 U15780 ( .A1(n13769), .A2(n13768), .ZN(n13953) );
  NAND3_X1 U15781 ( .A1(n13953), .A2(n13952), .A3(n15072), .ZN(n13770) );
  OAI211_X1 U15782 ( .C1(n13957), .C2(n15075), .A(n13771), .B(n13770), .ZN(
        P2_U3238) );
  XNOR2_X1 U15783 ( .A(n13772), .B(n13781), .ZN(n13774) );
  AOI21_X1 U15784 ( .B1(n13774), .B2(n13891), .A(n13773), .ZN(n13961) );
  INV_X1 U15785 ( .A(n13775), .ZN(n13776) );
  AOI211_X1 U15786 ( .C1(n13960), .C2(n13794), .A(n13777), .B(n13776), .ZN(
        n13959) );
  AOI22_X1 U15787 ( .A1(n13778), .A2(n15062), .B1(n15075), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n13779) );
  OAI21_X1 U15788 ( .B1(n13780), .B2(n15069), .A(n13779), .ZN(n13784) );
  XNOR2_X1 U15789 ( .A(n13782), .B(n13781), .ZN(n13963) );
  NOR2_X1 U15790 ( .A1(n13963), .A2(n13871), .ZN(n13783) );
  AOI211_X1 U15791 ( .C1(n13959), .C2(n15064), .A(n13784), .B(n13783), .ZN(
        n13785) );
  OAI21_X1 U15792 ( .B1(n15075), .B2(n13961), .A(n13785), .ZN(P2_U3239) );
  OR2_X1 U15793 ( .A1(n13786), .A2(n13791), .ZN(n13787) );
  NAND2_X1 U15794 ( .A1(n13788), .A2(n13787), .ZN(n13790) );
  AOI21_X1 U15795 ( .B1(n13790), .B2(n13891), .A(n13789), .ZN(n13968) );
  XNOR2_X1 U15796 ( .A(n13792), .B(n13791), .ZN(n13965) );
  NAND2_X1 U15797 ( .A1(n13809), .A2(n13964), .ZN(n13793) );
  NAND3_X1 U15798 ( .A1(n13794), .A2(n9326), .A3(n13793), .ZN(n13966) );
  INV_X1 U15799 ( .A(n13795), .ZN(n13796) );
  AOI22_X1 U15800 ( .A1(P2_REG2_REG_25__SCAN_IN), .A2(n15075), .B1(n13796), 
        .B2(n15062), .ZN(n13798) );
  NAND2_X1 U15801 ( .A1(n13964), .A2(n13927), .ZN(n13797) );
  OAI211_X1 U15802 ( .C1(n13966), .C2(n13866), .A(n13798), .B(n13797), .ZN(
        n13799) );
  AOI21_X1 U15803 ( .B1(n13965), .B2(n15072), .A(n13799), .ZN(n13800) );
  OAI21_X1 U15804 ( .B1(n13968), .B2(n15075), .A(n13800), .ZN(P2_U3240) );
  XNOR2_X1 U15805 ( .A(n13802), .B(n13801), .ZN(n13971) );
  NAND3_X1 U15806 ( .A1(n13818), .A2(n7199), .A3(n13803), .ZN(n13804) );
  AOI21_X1 U15807 ( .B1(n13805), .B2(n13804), .A(n13875), .ZN(n13806) );
  AOI211_X1 U15808 ( .C1(n13808), .C2(n13971), .A(n13807), .B(n13806), .ZN(
        n13975) );
  INV_X1 U15809 ( .A(n13809), .ZN(n13810) );
  AOI211_X1 U15810 ( .C1(n13973), .C2(n13830), .A(n6649), .B(n13810), .ZN(
        n13972) );
  NAND2_X1 U15811 ( .A1(n13972), .A2(n13923), .ZN(n13814) );
  INV_X1 U15812 ( .A(n13811), .ZN(n13812) );
  AOI22_X1 U15813 ( .A1(n15075), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13812), 
        .B2(n15062), .ZN(n13813) );
  OAI211_X1 U15814 ( .C1(n13815), .C2(n15069), .A(n13814), .B(n13813), .ZN(
        n13816) );
  AOI21_X1 U15815 ( .B1(n13925), .B2(n13971), .A(n13816), .ZN(n13817) );
  OAI21_X1 U15816 ( .B1(n13975), .B2(n15075), .A(n13817), .ZN(P2_U3241) );
  INV_X1 U15817 ( .A(n13818), .ZN(n13819) );
  AOI21_X1 U15818 ( .B1(n13820), .B2(n6484), .A(n13819), .ZN(n13822) );
  OAI21_X1 U15819 ( .B1(n13822), .B2(n13875), .A(n13821), .ZN(n13978) );
  NAND2_X1 U15820 ( .A1(n13978), .A2(n13868), .ZN(n13834) );
  NAND2_X1 U15821 ( .A1(n15075), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n13823) );
  OAI21_X1 U15822 ( .B1(n13825), .B2(n13824), .A(n13823), .ZN(n13826) );
  AOI21_X1 U15823 ( .B1(n13977), .B2(n13927), .A(n13826), .ZN(n13833) );
  XNOR2_X1 U15824 ( .A(n13828), .B(n13827), .ZN(n13980) );
  NAND2_X1 U15825 ( .A1(n13980), .A2(n15072), .ZN(n13832) );
  NAND2_X1 U15826 ( .A1(n13977), .A2(n13843), .ZN(n13829) );
  NAND2_X1 U15827 ( .A1(n13979), .A2(n13923), .ZN(n13831) );
  NAND4_X1 U15828 ( .A1(n13834), .A2(n13833), .A3(n13832), .A4(n13831), .ZN(
        P2_U3242) );
  XNOR2_X1 U15829 ( .A(n13835), .B(n13841), .ZN(n13837) );
  OAI21_X1 U15830 ( .B1(n13837), .B2(n13875), .A(n13836), .ZN(n13983) );
  INV_X1 U15831 ( .A(n13983), .ZN(n13853) );
  INV_X1 U15832 ( .A(n13838), .ZN(n13839) );
  AOI21_X1 U15833 ( .B1(n13841), .B2(n13840), .A(n13839), .ZN(n13985) );
  INV_X1 U15834 ( .A(n13842), .ZN(n13862) );
  INV_X1 U15835 ( .A(n13843), .ZN(n13844) );
  AOI211_X1 U15836 ( .C1(n13846), .C2(n13862), .A(n13845), .B(n13844), .ZN(
        n13984) );
  NAND2_X1 U15837 ( .A1(n13984), .A2(n13923), .ZN(n13850) );
  INV_X1 U15838 ( .A(n13847), .ZN(n13848) );
  AOI22_X1 U15839 ( .A1(n15075), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13848), 
        .B2(n15062), .ZN(n13849) );
  OAI211_X1 U15840 ( .C1(n14047), .C2(n15069), .A(n13850), .B(n13849), .ZN(
        n13851) );
  AOI21_X1 U15841 ( .B1(n13985), .B2(n15072), .A(n13851), .ZN(n13852) );
  OAI21_X1 U15842 ( .B1(n13853), .B2(n15075), .A(n13852), .ZN(P2_U3243) );
  XNOR2_X1 U15843 ( .A(n13854), .B(n13855), .ZN(n13990) );
  NAND2_X1 U15844 ( .A1(n13856), .A2(n13855), .ZN(n13857) );
  NAND3_X1 U15845 ( .A1(n13858), .A2(n13891), .A3(n13857), .ZN(n13860) );
  AND2_X1 U15846 ( .A1(n13860), .A2(n13859), .ZN(n13989) );
  INV_X1 U15847 ( .A(n13989), .ZN(n13869) );
  AOI21_X1 U15848 ( .B1(n13879), .B2(n14050), .A(n6649), .ZN(n13861) );
  NAND2_X1 U15849 ( .A1(n13862), .A2(n13861), .ZN(n13988) );
  AOI22_X1 U15850 ( .A1(n15075), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13863), 
        .B2(n15062), .ZN(n13865) );
  NAND2_X1 U15851 ( .A1(n14050), .A2(n13927), .ZN(n13864) );
  OAI211_X1 U15852 ( .C1(n13988), .C2(n13866), .A(n13865), .B(n13864), .ZN(
        n13867) );
  AOI21_X1 U15853 ( .B1(n13869), .B2(n13868), .A(n13867), .ZN(n13870) );
  OAI21_X1 U15854 ( .B1(n13871), .B2(n13990), .A(n13870), .ZN(P2_U3244) );
  XNOR2_X1 U15855 ( .A(n13873), .B(n13872), .ZN(n13876) );
  OAI21_X1 U15856 ( .B1(n13876), .B2(n13875), .A(n13874), .ZN(n13994) );
  INV_X1 U15857 ( .A(n13994), .ZN(n13888) );
  XNOR2_X1 U15858 ( .A(n13878), .B(n13877), .ZN(n13996) );
  INV_X1 U15859 ( .A(n13879), .ZN(n13880) );
  AOI211_X1 U15860 ( .C1(n13881), .C2(n13897), .A(n6649), .B(n13880), .ZN(
        n13995) );
  NAND2_X1 U15861 ( .A1(n13995), .A2(n13923), .ZN(n13885) );
  INV_X1 U15862 ( .A(n13882), .ZN(n13883) );
  AOI22_X1 U15863 ( .A1(n15075), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13883), 
        .B2(n15062), .ZN(n13884) );
  OAI211_X1 U15864 ( .C1(n6948), .C2(n15069), .A(n13885), .B(n13884), .ZN(
        n13886) );
  AOI21_X1 U15865 ( .B1(n15072), .B2(n13996), .A(n13886), .ZN(n13887) );
  OAI21_X1 U15866 ( .B1(n13888), .B2(n15075), .A(n13887), .ZN(P2_U3245) );
  OAI21_X1 U15867 ( .B1(n13890), .B2(n13896), .A(n13889), .ZN(n13892) );
  NAND2_X1 U15868 ( .A1(n13892), .A2(n13891), .ZN(n13894) );
  NAND2_X1 U15869 ( .A1(n13894), .A2(n13893), .ZN(n13999) );
  INV_X1 U15870 ( .A(n13999), .ZN(n13905) );
  AOI21_X1 U15871 ( .B1(n13896), .B2(n13895), .A(n6546), .ZN(n14001) );
  AOI211_X1 U15872 ( .C1(n13899), .C2(n13898), .A(n6649), .B(n6949), .ZN(
        n14000) );
  NAND2_X1 U15873 ( .A1(n14000), .A2(n13923), .ZN(n13902) );
  AOI22_X1 U15874 ( .A1(n15075), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13900), 
        .B2(n15062), .ZN(n13901) );
  OAI211_X1 U15875 ( .C1(n14059), .C2(n15069), .A(n13902), .B(n13901), .ZN(
        n13903) );
  AOI21_X1 U15876 ( .B1(n14001), .B2(n15072), .A(n13903), .ZN(n13904) );
  OAI21_X1 U15877 ( .B1(n13905), .B2(n15075), .A(n13904), .ZN(P2_U3246) );
  AOI22_X1 U15878 ( .A1(n15064), .A2(n13907), .B1(n15072), .B2(n13906), .ZN(
        n13913) );
  AOI22_X1 U15879 ( .A1(n13927), .A2(n13908), .B1(n15062), .B2(n9097), .ZN(
        n13912) );
  MUX2_X1 U15880 ( .A(n13910), .B(n13909), .S(n15075), .Z(n13911) );
  NAND3_X1 U15881 ( .A1(n13913), .A2(n13912), .A3(n13911), .ZN(P2_U3262) );
  AOI22_X1 U15882 ( .A1(n15064), .A2(n13915), .B1(n15072), .B2(n13914), .ZN(
        n13921) );
  AOI22_X1 U15883 ( .A1(n13927), .A2(n13916), .B1(n15062), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n13920) );
  MUX2_X1 U15884 ( .A(n13918), .B(n13917), .S(n15075), .Z(n13919) );
  NAND3_X1 U15885 ( .A1(n13921), .A2(n13920), .A3(n13919), .ZN(P2_U3263) );
  AOI22_X1 U15886 ( .A1(n13925), .A2(n13924), .B1(n13923), .B2(n13922), .ZN(
        n13932) );
  AOI22_X1 U15887 ( .A1(n13927), .A2(n13926), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n15062), .ZN(n13931) );
  MUX2_X1 U15888 ( .A(n13929), .B(n13928), .S(n15075), .Z(n13930) );
  NAND3_X1 U15889 ( .A1(n13932), .A2(n13931), .A3(n13930), .ZN(P2_U3264) );
  INV_X1 U15890 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13935) );
  NOR2_X1 U15891 ( .A1(n13934), .A2(n13933), .ZN(n14021) );
  MUX2_X1 U15892 ( .A(n13935), .B(n14021), .S(n15112), .Z(n13936) );
  OAI21_X1 U15893 ( .B1(n14024), .B2(n14015), .A(n13936), .ZN(P2_U3530) );
  INV_X1 U15894 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13939) );
  AND2_X1 U15895 ( .A1(n13938), .A2(n13937), .ZN(n14025) );
  MUX2_X1 U15896 ( .A(n13939), .B(n14025), .S(n15112), .Z(n13942) );
  NAND2_X1 U15897 ( .A1(n13940), .A2(n13992), .ZN(n13941) );
  NAND2_X1 U15898 ( .A1(n13942), .A2(n13941), .ZN(P2_U3529) );
  AOI21_X1 U15899 ( .B1(n15098), .B2(n13944), .A(n13943), .ZN(n13945) );
  MUX2_X1 U15900 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n14029), .S(n15112), .Z(
        P2_U3528) );
  OAI21_X1 U15901 ( .B1(n14032), .B2(n14015), .A(n13951), .ZN(P2_U3527) );
  NAND3_X1 U15902 ( .A1(n13953), .A2(n14012), .A3(n13952), .ZN(n13958) );
  NAND2_X1 U15903 ( .A1(n13954), .A2(n15098), .ZN(n13956) );
  NAND4_X1 U15904 ( .A1(n13958), .A2(n13957), .A3(n13956), .A4(n13955), .ZN(
        n14033) );
  MUX2_X1 U15905 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14033), .S(n15112), .Z(
        P2_U3526) );
  AOI21_X1 U15906 ( .B1(n15098), .B2(n13960), .A(n13959), .ZN(n13962) );
  OAI211_X1 U15907 ( .C1(n15093), .C2(n13963), .A(n13962), .B(n13961), .ZN(
        n14034) );
  MUX2_X1 U15908 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14034), .S(n15112), .Z(
        P2_U3525) );
  INV_X1 U15909 ( .A(n13964), .ZN(n14038) );
  NAND2_X1 U15910 ( .A1(n13965), .A2(n14012), .ZN(n13967) );
  AND3_X1 U15911 ( .A1(n13968), .A2(n13967), .A3(n13966), .ZN(n14035) );
  MUX2_X1 U15912 ( .A(n13969), .B(n14035), .S(n15112), .Z(n13970) );
  OAI21_X1 U15913 ( .B1(n14038), .B2(n14015), .A(n13970), .ZN(P2_U3524) );
  INV_X1 U15914 ( .A(n13971), .ZN(n13976) );
  AOI21_X1 U15915 ( .B1(n15098), .B2(n13973), .A(n13972), .ZN(n13974) );
  OAI211_X1 U15916 ( .C1(n13976), .C2(n15101), .A(n13975), .B(n13974), .ZN(
        n14039) );
  MUX2_X1 U15917 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14039), .S(n15112), .Z(
        P2_U3523) );
  INV_X1 U15918 ( .A(n13977), .ZN(n14043) );
  AOI211_X1 U15919 ( .C1(n13980), .C2(n14012), .A(n13979), .B(n13978), .ZN(
        n14040) );
  MUX2_X1 U15920 ( .A(n13981), .B(n14040), .S(n15112), .Z(n13982) );
  OAI21_X1 U15921 ( .B1(n14043), .B2(n14015), .A(n13982), .ZN(P2_U3522) );
  AOI211_X1 U15922 ( .C1(n13985), .C2(n14012), .A(n13984), .B(n13983), .ZN(
        n14044) );
  MUX2_X1 U15923 ( .A(n13986), .B(n14044), .S(n15112), .Z(n13987) );
  OAI21_X1 U15924 ( .B1(n14047), .B2(n14015), .A(n13987), .ZN(P2_U3521) );
  OAI211_X1 U15925 ( .C1(n15093), .C2(n13990), .A(n13989), .B(n13988), .ZN(
        n14048) );
  MUX2_X1 U15926 ( .A(n14048), .B(P2_REG1_REG_21__SCAN_IN), .S(n15109), .Z(
        n13991) );
  AOI21_X1 U15927 ( .B1(n13992), .B2(n14050), .A(n13991), .ZN(n13993) );
  INV_X1 U15928 ( .A(n13993), .ZN(P2_U3520) );
  AOI211_X1 U15929 ( .C1(n14012), .C2(n13996), .A(n13995), .B(n13994), .ZN(
        n14053) );
  MUX2_X1 U15930 ( .A(n13997), .B(n14053), .S(n15112), .Z(n13998) );
  OAI21_X1 U15931 ( .B1(n6948), .B2(n14015), .A(n13998), .ZN(P2_U3519) );
  AOI211_X1 U15932 ( .C1(n14001), .C2(n14012), .A(n14000), .B(n13999), .ZN(
        n14056) );
  MUX2_X1 U15933 ( .A(n14002), .B(n14056), .S(n15112), .Z(n14003) );
  OAI21_X1 U15934 ( .B1(n14059), .B2(n14015), .A(n14003), .ZN(P2_U3518) );
  AOI211_X1 U15935 ( .C1(n15098), .C2(n14006), .A(n14005), .B(n14004), .ZN(
        n14007) );
  OAI21_X1 U15936 ( .B1(n15093), .B2(n14008), .A(n14007), .ZN(n14060) );
  MUX2_X1 U15937 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14060), .S(n15112), .Z(
        P2_U3517) );
  AOI211_X1 U15938 ( .C1(n14012), .C2(n14011), .A(n14010), .B(n14009), .ZN(
        n14061) );
  MUX2_X1 U15939 ( .A(n14013), .B(n14061), .S(n15112), .Z(n14014) );
  OAI21_X1 U15940 ( .B1(n14065), .B2(n14015), .A(n14014), .ZN(P2_U3516) );
  AOI21_X1 U15941 ( .B1(n15098), .B2(n14017), .A(n14016), .ZN(n14018) );
  OAI211_X1 U15942 ( .C1(n15093), .C2(n14020), .A(n14019), .B(n14018), .ZN(
        n14066) );
  MUX2_X1 U15943 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n14066), .S(n15112), .Z(
        P2_U3512) );
  MUX2_X1 U15944 ( .A(n14022), .B(n14021), .S(n15106), .Z(n14023) );
  OAI21_X1 U15945 ( .B1(n14024), .B2(n14064), .A(n14023), .ZN(P2_U3498) );
  INV_X1 U15946 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14026) );
  MUX2_X1 U15947 ( .A(n14026), .B(n14025), .S(n15106), .Z(n14027) );
  OAI21_X1 U15948 ( .B1(n14028), .B2(n14064), .A(n14027), .ZN(P2_U3497) );
  MUX2_X1 U15949 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n14029), .S(n15106), .Z(
        P2_U3496) );
  INV_X1 U15950 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n14030) );
  OAI21_X1 U15951 ( .B1(n14032), .B2(n14064), .A(n14031), .ZN(P2_U3495) );
  MUX2_X1 U15952 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14033), .S(n15106), .Z(
        P2_U3494) );
  MUX2_X1 U15953 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14034), .S(n15106), .Z(
        P2_U3493) );
  INV_X1 U15954 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14036) );
  MUX2_X1 U15955 ( .A(n14036), .B(n14035), .S(n15106), .Z(n14037) );
  OAI21_X1 U15956 ( .B1(n14038), .B2(n14064), .A(n14037), .ZN(P2_U3492) );
  MUX2_X1 U15957 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14039), .S(n15106), .Z(
        P2_U3491) );
  INV_X1 U15958 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n14041) );
  MUX2_X1 U15959 ( .A(n14041), .B(n14040), .S(n15106), .Z(n14042) );
  OAI21_X1 U15960 ( .B1(n14043), .B2(n14064), .A(n14042), .ZN(P2_U3490) );
  INV_X1 U15961 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n14045) );
  MUX2_X1 U15962 ( .A(n14045), .B(n14044), .S(n15106), .Z(n14046) );
  OAI21_X1 U15963 ( .B1(n14047), .B2(n14064), .A(n14046), .ZN(P2_U3489) );
  MUX2_X1 U15964 ( .A(n14048), .B(P2_REG0_REG_21__SCAN_IN), .S(n15104), .Z(
        n14049) );
  AOI21_X1 U15965 ( .B1(n14051), .B2(n14050), .A(n14049), .ZN(n14052) );
  INV_X1 U15966 ( .A(n14052), .ZN(P2_U3488) );
  INV_X1 U15967 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n14054) );
  MUX2_X1 U15968 ( .A(n14054), .B(n14053), .S(n15106), .Z(n14055) );
  OAI21_X1 U15969 ( .B1(n6948), .B2(n14064), .A(n14055), .ZN(P2_U3487) );
  INV_X1 U15970 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14057) );
  MUX2_X1 U15971 ( .A(n14057), .B(n14056), .S(n15106), .Z(n14058) );
  OAI21_X1 U15972 ( .B1(n14059), .B2(n14064), .A(n14058), .ZN(P2_U3486) );
  MUX2_X1 U15973 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14060), .S(n15106), .Z(
        P2_U3484) );
  INV_X1 U15974 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14062) );
  MUX2_X1 U15975 ( .A(n14062), .B(n14061), .S(n15106), .Z(n14063) );
  OAI21_X1 U15976 ( .B1(n14065), .B2(n14064), .A(n14063), .ZN(P2_U3481) );
  MUX2_X1 U15977 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n14066), .S(n15106), .Z(
        P2_U3469) );
  INV_X1 U15978 ( .A(n14067), .ZN(n14680) );
  NOR4_X1 U15979 ( .A1(n8591), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14068), .A4(
        P2_U3088), .ZN(n14069) );
  AOI21_X1 U15980 ( .B1(n14070), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14069), 
        .ZN(n14071) );
  OAI21_X1 U15981 ( .B1(n14680), .B2(n14088), .A(n14071), .ZN(P2_U3296) );
  OAI222_X1 U15982 ( .A1(n14088), .A2(n14074), .B1(P2_U3088), .B2(n14073), 
        .C1(n14072), .C2(n14086), .ZN(P2_U3297) );
  OAI222_X1 U15983 ( .A1(n14088), .A2(n14077), .B1(P2_U3088), .B2(n14076), 
        .C1(n14075), .C2(n14086), .ZN(P2_U3298) );
  NAND2_X1 U15984 ( .A1(n11488), .A2(n14078), .ZN(n14080) );
  OAI211_X1 U15985 ( .C1(n14086), .C2(n14081), .A(n14080), .B(n14079), .ZN(
        P2_U3299) );
  INV_X1 U15986 ( .A(n14082), .ZN(n14687) );
  OAI222_X1 U15987 ( .A1(P2_U3088), .A2(n14084), .B1(n14086), .B2(n14083), 
        .C1(n14088), .C2(n14687), .ZN(P2_U3301) );
  INV_X1 U15988 ( .A(n14085), .ZN(n14695) );
  OAI222_X1 U15989 ( .A1(n14089), .A2(P2_U3088), .B1(n14088), .B2(n14695), 
        .C1(n14087), .C2(n14086), .ZN(P2_U3302) );
  INV_X1 U15990 ( .A(n14090), .ZN(n14091) );
  MUX2_X1 U15991 ( .A(n14091), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI211_X1 U15992 ( .C1(n14094), .C2(n14093), .A(n14092), .B(n14809), .ZN(
        n14101) );
  AOI22_X1 U15993 ( .A1(n14217), .A2(n14259), .B1(P1_REG3_REG_7__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14100) );
  INV_X1 U15994 ( .A(n14095), .ZN(n14097) );
  AOI22_X1 U15995 ( .A1(n14236), .A2(n14097), .B1(n14879), .B2(n14096), .ZN(
        n14099) );
  NAND2_X1 U15996 ( .A1(n14115), .A2(n14261), .ZN(n14098) );
  NAND4_X1 U15997 ( .A1(n14101), .A2(n14100), .A3(n14099), .A4(n14098), .ZN(
        P1_U3213) );
  OAI22_X1 U15998 ( .A1(n14870), .A2(n14103), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14102), .ZN(n14104) );
  AOI21_X1 U15999 ( .B1(n14217), .B2(n14345), .A(n14104), .ZN(n14105) );
  OAI21_X1 U16000 ( .B1(n14883), .B2(n14350), .A(n14105), .ZN(n14106) );
  AOI21_X1 U16001 ( .B1(n14572), .B2(n14879), .A(n14106), .ZN(n14107) );
  OAI21_X1 U16002 ( .B1(n14108), .B2(n14875), .A(n14107), .ZN(P1_U3214) );
  AOI21_X1 U16003 ( .B1(n14111), .B2(n14110), .A(n14109), .ZN(n14121) );
  OAI22_X1 U16004 ( .A1(n14871), .A2(n14113), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14112), .ZN(n14114) );
  AOI21_X1 U16005 ( .B1(n14115), .B2(n14254), .A(n14114), .ZN(n14116) );
  OAI21_X1 U16006 ( .B1(n14883), .B2(n14117), .A(n14116), .ZN(n14118) );
  AOI21_X1 U16007 ( .B1(n14119), .B2(n14879), .A(n14118), .ZN(n14120) );
  OAI21_X1 U16008 ( .B1(n14121), .B2(n14875), .A(n14120), .ZN(P1_U3215) );
  XOR2_X1 U16009 ( .A(n14123), .B(n14122), .Z(n14129) );
  AND2_X1 U16010 ( .A1(n14420), .A2(n14961), .ZN(n14600) );
  OR2_X1 U16011 ( .A1(n14150), .A2(n14517), .ZN(n14125) );
  NAND2_X1 U16012 ( .A1(n14244), .A2(n14921), .ZN(n14124) );
  NAND2_X1 U16013 ( .A1(n14125), .A2(n14124), .ZN(n14598) );
  AOI22_X1 U16014 ( .A1(n14225), .A2(n14598), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14126) );
  OAI21_X1 U16015 ( .B1(n14883), .B2(n14421), .A(n14126), .ZN(n14127) );
  AOI21_X1 U16016 ( .B1(n14600), .B2(n14815), .A(n14127), .ZN(n14128) );
  OAI21_X1 U16017 ( .B1(n14129), .B2(n14875), .A(n14128), .ZN(P1_U3216) );
  AOI21_X1 U16018 ( .B1(n14131), .B2(n14130), .A(n14875), .ZN(n14133) );
  NAND2_X1 U16019 ( .A1(n14133), .A2(n14132), .ZN(n14139) );
  AOI22_X1 U16020 ( .A1(n14879), .A2(n14135), .B1(n14225), .B2(n14134), .ZN(
        n14138) );
  MUX2_X1 U16021 ( .A(P1_STATE_REG_SCAN_IN), .B(n14883), .S(n14136), .Z(n14137) );
  NAND3_X1 U16022 ( .A1(n14139), .A2(n14138), .A3(n14137), .ZN(P1_U3218) );
  INV_X1 U16023 ( .A(n14489), .ZN(n14626) );
  OAI211_X1 U16024 ( .C1(n14142), .C2(n14141), .A(n14140), .B(n14809), .ZN(
        n14145) );
  AOI22_X1 U16025 ( .A1(n14247), .A2(n14921), .B1(n14394), .B2(n14249), .ZN(
        n14624) );
  NAND2_X1 U16026 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14328)
         );
  OAI21_X1 U16027 ( .B1(n14624), .B2(n14233), .A(n14328), .ZN(n14143) );
  AOI21_X1 U16028 ( .B1(n14481), .B2(n14236), .A(n14143), .ZN(n14144) );
  OAI211_X1 U16029 ( .C1(n14626), .C2(n14239), .A(n14145), .B(n14144), .ZN(
        P1_U3219) );
  INV_X1 U16030 ( .A(n14146), .ZN(n14147) );
  AOI21_X1 U16031 ( .B1(n14149), .B2(n14148), .A(n14147), .ZN(n14156) );
  NOR2_X1 U16032 ( .A1(n14883), .A2(n14448), .ZN(n14154) );
  NOR2_X1 U16033 ( .A1(n14150), .A2(n14637), .ZN(n14151) );
  AOI21_X1 U16034 ( .B1(n14247), .B2(n14394), .A(n14151), .ZN(n14442) );
  INV_X1 U16035 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14152) );
  OAI22_X1 U16036 ( .A1(n14442), .A2(n14233), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14152), .ZN(n14153) );
  AOI211_X1 U16037 ( .C1(n14451), .C2(n14879), .A(n14154), .B(n14153), .ZN(
        n14155) );
  OAI21_X1 U16038 ( .B1(n14156), .B2(n14875), .A(n14155), .ZN(P1_U3223) );
  XOR2_X1 U16039 ( .A(n14158), .B(n14157), .Z(n14164) );
  NAND2_X1 U16040 ( .A1(n14244), .A2(n14394), .ZN(n14160) );
  NAND2_X1 U16041 ( .A1(n14346), .A2(n14921), .ZN(n14159) );
  NAND2_X1 U16042 ( .A1(n14160), .A2(n14159), .ZN(n14585) );
  AOI22_X1 U16043 ( .A1(n14225), .A2(n14585), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14161) );
  OAI21_X1 U16044 ( .B1(n14883), .B2(n14376), .A(n14161), .ZN(n14162) );
  AOI21_X1 U16045 ( .B1(n14586), .B2(n14879), .A(n14162), .ZN(n14163) );
  OAI21_X1 U16046 ( .B1(n14164), .B2(n14875), .A(n14163), .ZN(P1_U3225) );
  INV_X1 U16047 ( .A(n14165), .ZN(n14166) );
  AOI21_X1 U16048 ( .B1(n14168), .B2(n14167), .A(n14166), .ZN(n14175) );
  AOI22_X1 U16049 ( .A1(n14225), .A2(n14169), .B1(P1_REG3_REG_16__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14170) );
  OAI21_X1 U16050 ( .B1(n14883), .B2(n14171), .A(n14170), .ZN(n14172) );
  AOI21_X1 U16051 ( .B1(n14173), .B2(n14879), .A(n14172), .ZN(n14174) );
  OAI21_X1 U16052 ( .B1(n14175), .B2(n14875), .A(n14174), .ZN(P1_U3226) );
  XOR2_X1 U16053 ( .A(n14177), .B(n14176), .Z(n14183) );
  NOR2_X1 U16054 ( .A1(n14883), .A2(n14522), .ZN(n14181) );
  NAND2_X1 U16055 ( .A1(n14217), .A2(n14249), .ZN(n14179) );
  NAND2_X1 U16056 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14293)
         );
  OAI211_X1 U16057 ( .C1(n14518), .C2(n14870), .A(n14179), .B(n14293), .ZN(
        n14180) );
  AOI211_X1 U16058 ( .C1(n14636), .C2(n14879), .A(n14181), .B(n14180), .ZN(
        n14182) );
  OAI21_X1 U16059 ( .B1(n14183), .B2(n14875), .A(n14182), .ZN(P1_U3228) );
  INV_X1 U16060 ( .A(n14815), .ZN(n14193) );
  NAND2_X1 U16061 ( .A1(n14403), .A2(n14961), .ZN(n14592) );
  XNOR2_X1 U16062 ( .A(n14185), .B(n14184), .ZN(n14186) );
  NAND2_X1 U16063 ( .A1(n14186), .A2(n14809), .ZN(n14192) );
  OAI22_X1 U16064 ( .A1(n14870), .A2(n14188), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14187), .ZN(n14190) );
  NOR2_X1 U16065 ( .A1(n14883), .A2(n14401), .ZN(n14189) );
  AOI211_X1 U16066 ( .C1(n14217), .C2(n14392), .A(n14190), .B(n14189), .ZN(
        n14191) );
  OAI211_X1 U16067 ( .C1(n14193), .C2(n14592), .A(n14192), .B(n14191), .ZN(
        P1_U3229) );
  INV_X1 U16068 ( .A(n14470), .ZN(n14618) );
  OAI211_X1 U16069 ( .C1(n14196), .C2(n14195), .A(n14194), .B(n14809), .ZN(
        n14201) );
  AND2_X1 U16070 ( .A1(n14246), .A2(n14921), .ZN(n14197) );
  AOI21_X1 U16071 ( .B1(n14248), .B2(n14394), .A(n14197), .ZN(n14617) );
  OAI22_X1 U16072 ( .A1(n14617), .A2(n14233), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14198), .ZN(n14199) );
  AOI21_X1 U16073 ( .B1(n14466), .B2(n14236), .A(n14199), .ZN(n14200) );
  OAI211_X1 U16074 ( .C1(n14618), .C2(n14239), .A(n14201), .B(n14200), .ZN(
        P1_U3233) );
  OAI21_X1 U16075 ( .B1(n14204), .B2(n14203), .A(n14202), .ZN(n14205) );
  NAND2_X1 U16076 ( .A1(n14205), .A2(n14809), .ZN(n14212) );
  INV_X1 U16077 ( .A(n14433), .ZN(n14210) );
  NAND2_X1 U16078 ( .A1(n14246), .A2(n14394), .ZN(n14207) );
  NAND2_X1 U16079 ( .A1(n14393), .A2(n14921), .ZN(n14206) );
  AND2_X1 U16080 ( .A1(n14207), .A2(n14206), .ZN(n14604) );
  INV_X1 U16081 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14208) );
  OAI22_X1 U16082 ( .A1(n14233), .A2(n14604), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14208), .ZN(n14209) );
  AOI21_X1 U16083 ( .B1(n14236), .B2(n14210), .A(n14209), .ZN(n14211) );
  OAI211_X1 U16084 ( .C1(n14239), .C2(n14606), .A(n14212), .B(n14211), .ZN(
        P1_U3235) );
  XOR2_X1 U16085 ( .A(n14214), .B(n14213), .Z(n14221) );
  OAI21_X1 U16086 ( .B1(n14870), .B2(n14493), .A(n14215), .ZN(n14216) );
  AOI21_X1 U16087 ( .B1(n14217), .B2(n14248), .A(n14216), .ZN(n14218) );
  OAI21_X1 U16088 ( .B1(n14883), .B2(n14503), .A(n14218), .ZN(n14219) );
  AOI21_X1 U16089 ( .B1(n14632), .B2(n14879), .A(n14219), .ZN(n14220) );
  OAI21_X1 U16090 ( .B1(n14221), .B2(n14875), .A(n14220), .ZN(P1_U3238) );
  NAND2_X1 U16091 ( .A1(n14392), .A2(n14394), .ZN(n14224) );
  NAND2_X1 U16092 ( .A1(n14243), .A2(n14921), .ZN(n14223) );
  NAND2_X1 U16093 ( .A1(n14224), .A2(n14223), .ZN(n14577) );
  AOI22_X1 U16094 ( .A1(n14225), .A2(n14577), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14226) );
  OAI21_X1 U16095 ( .B1(n14883), .B2(n14363), .A(n14226), .ZN(n14227) );
  AOI21_X1 U16096 ( .B1(n14578), .B2(n14879), .A(n14227), .ZN(n14228) );
  OAI21_X1 U16097 ( .B1(n14229), .B2(n14875), .A(n14228), .ZN(P1_U3240) );
  OAI211_X1 U16098 ( .C1(n14232), .C2(n14231), .A(n14230), .B(n14809), .ZN(
        n14238) );
  INV_X1 U16099 ( .A(n14542), .ZN(n14235) );
  AOI22_X1 U16100 ( .A1(n14394), .A2(n14253), .B1(n14251), .B2(n14921), .ZN(
        n14536) );
  NAND2_X1 U16101 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14909)
         );
  OAI21_X1 U16102 ( .B1(n14233), .B2(n14536), .A(n14909), .ZN(n14234) );
  AOI21_X1 U16103 ( .B1(n14236), .B2(n14235), .A(n14234), .ZN(n14237) );
  OAI211_X1 U16104 ( .C1(n14240), .C2(n14239), .A(n14238), .B(n14237), .ZN(
        P1_U3241) );
  MUX2_X1 U16105 ( .A(n14334), .B(P1_DATAO_REG_31__SCAN_IN), .S(n14266), .Z(
        P1_U3591) );
  MUX2_X1 U16106 ( .A(n14241), .B(P1_DATAO_REG_30__SCAN_IN), .S(n14266), .Z(
        P1_U3590) );
  MUX2_X1 U16107 ( .A(n14242), .B(P1_DATAO_REG_29__SCAN_IN), .S(n14266), .Z(
        P1_U3589) );
  MUX2_X1 U16108 ( .A(n14345), .B(P1_DATAO_REG_28__SCAN_IN), .S(n14266), .Z(
        P1_U3588) );
  MUX2_X1 U16109 ( .A(n14243), .B(P1_DATAO_REG_27__SCAN_IN), .S(n14266), .Z(
        P1_U3587) );
  MUX2_X1 U16110 ( .A(n14346), .B(P1_DATAO_REG_26__SCAN_IN), .S(n14266), .Z(
        P1_U3586) );
  MUX2_X1 U16111 ( .A(n14392), .B(P1_DATAO_REG_25__SCAN_IN), .S(n14266), .Z(
        P1_U3585) );
  MUX2_X1 U16112 ( .A(n14244), .B(P1_DATAO_REG_24__SCAN_IN), .S(n14266), .Z(
        P1_U3584) );
  MUX2_X1 U16113 ( .A(n14393), .B(P1_DATAO_REG_23__SCAN_IN), .S(n14266), .Z(
        P1_U3583) );
  MUX2_X1 U16114 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14245), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16115 ( .A(n14246), .B(P1_DATAO_REG_21__SCAN_IN), .S(n14266), .Z(
        P1_U3581) );
  MUX2_X1 U16116 ( .A(n14247), .B(P1_DATAO_REG_20__SCAN_IN), .S(n14266), .Z(
        P1_U3580) );
  MUX2_X1 U16117 ( .A(n14248), .B(P1_DATAO_REG_19__SCAN_IN), .S(n14266), .Z(
        P1_U3579) );
  MUX2_X1 U16118 ( .A(n14249), .B(P1_DATAO_REG_18__SCAN_IN), .S(n14266), .Z(
        P1_U3578) );
  MUX2_X1 U16119 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14250), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16120 ( .A(n14251), .B(P1_DATAO_REG_16__SCAN_IN), .S(n14266), .Z(
        P1_U3576) );
  MUX2_X1 U16121 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14252), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16122 ( .A(n14253), .B(P1_DATAO_REG_14__SCAN_IN), .S(n14266), .Z(
        P1_U3574) );
  MUX2_X1 U16123 ( .A(n14254), .B(P1_DATAO_REG_13__SCAN_IN), .S(n14266), .Z(
        P1_U3573) );
  MUX2_X1 U16124 ( .A(n14255), .B(P1_DATAO_REG_12__SCAN_IN), .S(n14266), .Z(
        P1_U3572) );
  MUX2_X1 U16125 ( .A(n14256), .B(P1_DATAO_REG_11__SCAN_IN), .S(n14266), .Z(
        P1_U3571) );
  MUX2_X1 U16126 ( .A(n14257), .B(P1_DATAO_REG_10__SCAN_IN), .S(n14266), .Z(
        P1_U3570) );
  MUX2_X1 U16127 ( .A(n14258), .B(P1_DATAO_REG_9__SCAN_IN), .S(n14266), .Z(
        P1_U3569) );
  MUX2_X1 U16128 ( .A(n14259), .B(P1_DATAO_REG_8__SCAN_IN), .S(n14266), .Z(
        P1_U3568) );
  MUX2_X1 U16129 ( .A(n14260), .B(P1_DATAO_REG_7__SCAN_IN), .S(n14266), .Z(
        P1_U3567) );
  MUX2_X1 U16130 ( .A(n14261), .B(P1_DATAO_REG_6__SCAN_IN), .S(n14266), .Z(
        P1_U3566) );
  MUX2_X1 U16131 ( .A(n14262), .B(P1_DATAO_REG_5__SCAN_IN), .S(n14266), .Z(
        P1_U3565) );
  MUX2_X1 U16132 ( .A(n14263), .B(P1_DATAO_REG_4__SCAN_IN), .S(n14266), .Z(
        P1_U3564) );
  MUX2_X1 U16133 ( .A(n14264), .B(P1_DATAO_REG_3__SCAN_IN), .S(n14266), .Z(
        P1_U3563) );
  MUX2_X1 U16134 ( .A(n9387), .B(P1_DATAO_REG_2__SCAN_IN), .S(n14266), .Z(
        P1_U3562) );
  MUX2_X1 U16135 ( .A(n6688), .B(P1_DATAO_REG_1__SCAN_IN), .S(n14266), .Z(
        P1_U3561) );
  MUX2_X1 U16136 ( .A(n14267), .B(P1_DATAO_REG_0__SCAN_IN), .S(n14266), .Z(
        P1_U3560) );
  OAI211_X1 U16137 ( .C1(n14270), .C2(n14269), .A(n14901), .B(n14268), .ZN(
        n14279) );
  OAI211_X1 U16138 ( .C1(n14273), .C2(n14272), .A(n14318), .B(n14271), .ZN(
        n14278) );
  AOI22_X1 U16139 ( .A1(n14891), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14277) );
  INV_X1 U16140 ( .A(n14274), .ZN(n14275) );
  NAND2_X1 U16141 ( .A1(n14903), .A2(n14275), .ZN(n14276) );
  NAND4_X1 U16142 ( .A1(n14279), .A2(n14278), .A3(n14277), .A4(n14276), .ZN(
        P1_U3244) );
  AND2_X1 U16143 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n14281) );
  NOR2_X1 U16144 ( .A1(n14320), .A2(n6865), .ZN(n14280) );
  AOI211_X1 U16145 ( .C1(n14891), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n14281), .B(
        n14280), .ZN(n14292) );
  OAI211_X1 U16146 ( .C1(n14284), .C2(n14283), .A(n14901), .B(n14282), .ZN(
        n14291) );
  OR3_X1 U16147 ( .A1(n14287), .A2(n14286), .A3(n14285), .ZN(n14288) );
  NAND3_X1 U16148 ( .A1(n14318), .A2(n14289), .A3(n14288), .ZN(n14290) );
  NAND3_X1 U16149 ( .A1(n14292), .A2(n14291), .A3(n14290), .ZN(P1_U3246) );
  OAI21_X1 U16150 ( .B1(n14911), .B2(n7462), .A(n14293), .ZN(n14294) );
  AOI21_X1 U16151 ( .B1(n14295), .B2(n14903), .A(n14294), .ZN(n14306) );
  OAI211_X1 U16152 ( .C1(n14298), .C2(n14297), .A(n14901), .B(n14296), .ZN(
        n14305) );
  NAND2_X1 U16153 ( .A1(n14300), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14299) );
  OAI21_X1 U16154 ( .B1(n14300), .B2(P1_REG2_REG_17__SCAN_IN), .A(n14299), 
        .ZN(n14302) );
  OAI211_X1 U16155 ( .C1(n14303), .C2(n14302), .A(n14318), .B(n14301), .ZN(
        n14304) );
  NAND3_X1 U16156 ( .A1(n14306), .A2(n14305), .A3(n14304), .ZN(P1_U3260) );
  NOR2_X1 U16157 ( .A1(n14308), .A2(n14307), .ZN(n14310) );
  NOR2_X1 U16158 ( .A1(n14310), .A2(n14309), .ZN(n14312) );
  XNOR2_X1 U16159 ( .A(n14312), .B(n14311), .ZN(n14324) );
  INV_X1 U16160 ( .A(n14324), .ZN(n14321) );
  NAND2_X1 U16161 ( .A1(n14314), .A2(n14313), .ZN(n14315) );
  NAND2_X1 U16162 ( .A1(n14316), .A2(n14315), .ZN(n14317) );
  XNOR2_X1 U16163 ( .A(n14317), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n14322) );
  NAND2_X1 U16164 ( .A1(n14322), .A2(n14318), .ZN(n14319) );
  OAI211_X1 U16165 ( .C1(n14321), .C2(n14323), .A(n14320), .B(n14319), .ZN(
        n14326) );
  OAI22_X1 U16166 ( .A1(n14324), .A2(n14323), .B1(n14322), .B2(n14906), .ZN(
        n14325) );
  MUX2_X1 U16167 ( .A(n14326), .B(n14325), .S(n14540), .Z(n14327) );
  INV_X1 U16168 ( .A(n14327), .ZN(n14329) );
  OAI211_X1 U16169 ( .C1(n7316), .C2(n14911), .A(n14329), .B(n14328), .ZN(
        P1_U3262) );
  XNOR2_X1 U16170 ( .A(n14552), .B(n14337), .ZN(n14332) );
  NAND2_X1 U16171 ( .A1(n14332), .A2(n14736), .ZN(n14551) );
  NAND2_X1 U16172 ( .A1(n14334), .A2(n14333), .ZN(n14553) );
  NOR2_X1 U16173 ( .A1(n14743), .A2(n14553), .ZN(n14340) );
  NOR2_X1 U16174 ( .A1(n14552), .A2(n14506), .ZN(n14335) );
  AOI211_X1 U16175 ( .C1(n14743), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14340), 
        .B(n14335), .ZN(n14336) );
  OAI21_X1 U16176 ( .B1(n14551), .B2(n14486), .A(n14336), .ZN(P1_U3263) );
  OAI211_X1 U16177 ( .C1(n14555), .C2(n14338), .A(n14337), .B(n14736), .ZN(
        n14554) );
  NOR2_X1 U16178 ( .A1(n14555), .A2(n14506), .ZN(n14339) );
  AOI211_X1 U16179 ( .C1(n14743), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14340), 
        .B(n14339), .ZN(n14341) );
  OAI21_X1 U16180 ( .B1(n14486), .B2(n14554), .A(n14341), .ZN(P1_U3264) );
  INV_X1 U16181 ( .A(n14575), .ZN(n14354) );
  AOI22_X1 U16182 ( .A1(n14394), .A2(n14346), .B1(n14345), .B2(n14921), .ZN(
        n14347) );
  AOI211_X1 U16183 ( .C1(n14572), .C2(n14361), .A(n14924), .B(n14348), .ZN(
        n14571) );
  NOR2_X1 U16184 ( .A1(n14349), .A2(n14506), .ZN(n14353) );
  OAI22_X1 U16185 ( .A1(n14544), .A2(n14351), .B1(n14350), .B2(n14541), .ZN(
        n14352) );
  AOI211_X1 U16186 ( .C1(n14571), .C2(n14739), .A(n14353), .B(n14352), .ZN(
        n14356) );
  NAND2_X1 U16187 ( .A1(n14354), .A2(n14740), .ZN(n14355) );
  OAI211_X1 U16188 ( .C1(n14574), .C2(n14743), .A(n14356), .B(n14355), .ZN(
        P1_U3266) );
  XNOR2_X1 U16189 ( .A(n14357), .B(n14359), .ZN(n14582) );
  OAI21_X1 U16190 ( .B1(n14360), .B2(n14359), .A(n14358), .ZN(n14579) );
  INV_X1 U16191 ( .A(n14361), .ZN(n14362) );
  AOI211_X1 U16192 ( .C1(n14578), .C2(n14374), .A(n14924), .B(n14362), .ZN(
        n14576) );
  AOI21_X1 U16193 ( .B1(n14576), .B2(n14540), .A(n14577), .ZN(n14367) );
  INV_X1 U16194 ( .A(n14363), .ZN(n14364) );
  AOI22_X1 U16195 ( .A1(n14743), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n14364), 
        .B2(n14732), .ZN(n14366) );
  NAND2_X1 U16196 ( .A1(n14578), .A2(n14733), .ZN(n14365) );
  OAI211_X1 U16197 ( .C1(n14367), .C2(n14743), .A(n14366), .B(n14365), .ZN(
        n14368) );
  AOI21_X1 U16198 ( .B1(n14480), .B2(n14579), .A(n14368), .ZN(n14369) );
  OAI21_X1 U16199 ( .B1(n14546), .B2(n14582), .A(n14369), .ZN(P1_U3267) );
  XNOR2_X1 U16200 ( .A(n14370), .B(n14373), .ZN(n14589) );
  AOI21_X1 U16201 ( .B1(n14373), .B2(n14372), .A(n14371), .ZN(n14583) );
  NAND2_X1 U16202 ( .A1(n14583), .A2(n14474), .ZN(n14384) );
  AOI21_X1 U16203 ( .B1(n14400), .B2(n14586), .A(n14924), .ZN(n14375) );
  AND2_X1 U16204 ( .A1(n14375), .A2(n14374), .ZN(n14584) );
  NAND2_X1 U16205 ( .A1(n14586), .A2(n14733), .ZN(n14381) );
  INV_X1 U16206 ( .A(n14585), .ZN(n14377) );
  OAI22_X1 U16207 ( .A1(n14743), .A2(n14377), .B1(n14376), .B2(n14541), .ZN(
        n14378) );
  INV_X1 U16208 ( .A(n14378), .ZN(n14380) );
  NAND2_X1 U16209 ( .A1(n14743), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n14379) );
  NAND3_X1 U16210 ( .A1(n14381), .A2(n14380), .A3(n14379), .ZN(n14382) );
  AOI21_X1 U16211 ( .B1(n14584), .B2(n14739), .A(n14382), .ZN(n14383) );
  OAI211_X1 U16212 ( .C1(n14589), .C2(n14476), .A(n14384), .B(n14383), .ZN(
        P1_U3268) );
  OAI211_X1 U16213 ( .C1(n14387), .C2(n14386), .A(n14385), .B(n14832), .ZN(
        n14397) );
  OR2_X1 U16214 ( .A1(n14389), .A2(n14388), .ZN(n14390) );
  NAND2_X1 U16215 ( .A1(n14391), .A2(n14390), .ZN(n14590) );
  NAND2_X1 U16216 ( .A1(n14590), .A2(n14729), .ZN(n14396) );
  AOI22_X1 U16217 ( .A1(n14394), .A2(n14393), .B1(n14392), .B2(n14921), .ZN(
        n14395) );
  NAND3_X1 U16218 ( .A1(n14397), .A2(n14396), .A3(n14395), .ZN(n14595) );
  INV_X1 U16219 ( .A(n14595), .ZN(n14408) );
  INV_X1 U16220 ( .A(n14419), .ZN(n14398) );
  AOI21_X1 U16221 ( .B1(n14403), .B2(n14398), .A(n14924), .ZN(n14399) );
  NAND2_X1 U16222 ( .A1(n14400), .A2(n14399), .ZN(n14591) );
  INV_X1 U16223 ( .A(n14401), .ZN(n14402) );
  AOI22_X1 U16224 ( .A1(n14743), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14402), 
        .B2(n14732), .ZN(n14405) );
  NAND2_X1 U16225 ( .A1(n14403), .A2(n14733), .ZN(n14404) );
  OAI211_X1 U16226 ( .C1(n14591), .C2(n14486), .A(n14405), .B(n14404), .ZN(
        n14406) );
  AOI21_X1 U16227 ( .B1(n14590), .B2(n14740), .A(n14406), .ZN(n14407) );
  OAI21_X1 U16228 ( .B1(n14408), .B2(n14743), .A(n14407), .ZN(P1_U3269) );
  OAI21_X1 U16229 ( .B1(n14411), .B2(n14410), .A(n14409), .ZN(n14412) );
  INV_X1 U16230 ( .A(n14412), .ZN(n14603) );
  OAI21_X1 U16231 ( .B1(n14415), .B2(n14414), .A(n14413), .ZN(n14416) );
  AND2_X1 U16232 ( .A1(n14416), .A2(n14832), .ZN(n14601) );
  OAI21_X1 U16233 ( .B1(n14601), .B2(n14598), .A(n14544), .ZN(n14427) );
  NAND2_X1 U16234 ( .A1(n14420), .A2(n14432), .ZN(n14417) );
  NAND2_X1 U16235 ( .A1(n14417), .A2(n14736), .ZN(n14418) );
  NOR2_X1 U16236 ( .A1(n14419), .A2(n14418), .ZN(n14599) );
  INV_X1 U16237 ( .A(n14420), .ZN(n14424) );
  INV_X1 U16238 ( .A(n14421), .ZN(n14422) );
  AOI22_X1 U16239 ( .A1(n14743), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n14422), 
        .B2(n14732), .ZN(n14423) );
  OAI21_X1 U16240 ( .B1(n14424), .B2(n14506), .A(n14423), .ZN(n14425) );
  AOI21_X1 U16241 ( .B1(n14599), .B2(n14739), .A(n14425), .ZN(n14426) );
  OAI211_X1 U16242 ( .C1(n14603), .C2(n14546), .A(n14427), .B(n14426), .ZN(
        P1_U3270) );
  XOR2_X1 U16243 ( .A(n14430), .B(n14428), .Z(n14610) );
  OAI21_X1 U16244 ( .B1(n14431), .B2(n14430), .A(n14429), .ZN(n14608) );
  OAI211_X1 U16245 ( .C1(n14606), .C2(n14447), .A(n14736), .B(n14432), .ZN(
        n14605) );
  OAI22_X1 U16246 ( .A1(n14743), .A2(n14604), .B1(n14433), .B2(n14541), .ZN(
        n14435) );
  NOR2_X1 U16247 ( .A1(n14606), .A2(n14506), .ZN(n14434) );
  AOI211_X1 U16248 ( .C1(n14743), .C2(P1_REG2_REG_22__SCAN_IN), .A(n14435), 
        .B(n14434), .ZN(n14436) );
  OAI21_X1 U16249 ( .B1(n14486), .B2(n14605), .A(n14436), .ZN(n14437) );
  AOI21_X1 U16250 ( .B1(n14608), .B2(n14474), .A(n14437), .ZN(n14438) );
  OAI21_X1 U16251 ( .B1(n14610), .B2(n14476), .A(n14438), .ZN(P1_U3271) );
  XNOR2_X1 U16252 ( .A(n14440), .B(n14439), .ZN(n14441) );
  NAND2_X1 U16253 ( .A1(n14441), .A2(n14832), .ZN(n14443) );
  NAND2_X1 U16254 ( .A1(n14443), .A2(n14442), .ZN(n14616) );
  INV_X1 U16255 ( .A(n14616), .ZN(n14455) );
  XNOR2_X1 U16256 ( .A(n14445), .B(n14444), .ZN(n14611) );
  OAI21_X1 U16257 ( .B1(n14465), .B2(n14614), .A(n14736), .ZN(n14446) );
  OR2_X1 U16258 ( .A1(n14447), .A2(n14446), .ZN(n14612) );
  OAI22_X1 U16259 ( .A1(n14544), .A2(n14449), .B1(n14448), .B2(n14541), .ZN(
        n14450) );
  AOI21_X1 U16260 ( .B1(n14451), .B2(n14733), .A(n14450), .ZN(n14452) );
  OAI21_X1 U16261 ( .B1(n14612), .B2(n14486), .A(n14452), .ZN(n14453) );
  AOI21_X1 U16262 ( .B1(n14611), .B2(n14474), .A(n14453), .ZN(n14454) );
  OAI21_X1 U16263 ( .B1(n14455), .B2(n14743), .A(n14454), .ZN(P1_U3272) );
  OAI21_X1 U16264 ( .B1(n14461), .B2(n14457), .A(n14456), .ZN(n14623) );
  INV_X1 U16265 ( .A(n14458), .ZN(n14459) );
  AOI21_X1 U16266 ( .B1(n14461), .B2(n14460), .A(n14459), .ZN(n14621) );
  NAND2_X1 U16267 ( .A1(n14462), .A2(n14470), .ZN(n14463) );
  NAND2_X1 U16268 ( .A1(n14463), .A2(n14736), .ZN(n14464) );
  NOR2_X1 U16269 ( .A1(n14465), .A2(n14464), .ZN(n14620) );
  NAND2_X1 U16270 ( .A1(n14620), .A2(n14739), .ZN(n14472) );
  NAND2_X1 U16271 ( .A1(n14466), .A2(n14732), .ZN(n14468) );
  NAND2_X1 U16272 ( .A1(n14743), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n14467) );
  OAI211_X1 U16273 ( .C1(n14617), .C2(n14743), .A(n14468), .B(n14467), .ZN(
        n14469) );
  AOI21_X1 U16274 ( .B1(n14470), .B2(n14733), .A(n14469), .ZN(n14471) );
  NAND2_X1 U16275 ( .A1(n14472), .A2(n14471), .ZN(n14473) );
  AOI21_X1 U16276 ( .B1(n14621), .B2(n14474), .A(n14473), .ZN(n14475) );
  OAI21_X1 U16277 ( .B1(n14476), .B2(n14623), .A(n14475), .ZN(P1_U3273) );
  XNOR2_X1 U16278 ( .A(n14477), .B(n14478), .ZN(n14630) );
  XNOR2_X1 U16279 ( .A(n14479), .B(n14478), .ZN(n14628) );
  NAND2_X1 U16280 ( .A1(n14628), .A2(n14480), .ZN(n14491) );
  INV_X1 U16281 ( .A(n14624), .ZN(n14482) );
  AOI22_X1 U16282 ( .A1(n14482), .A2(n14544), .B1(n14481), .B2(n14732), .ZN(
        n14483) );
  OAI21_X1 U16283 ( .B1(n14484), .B2(n14544), .A(n14483), .ZN(n14488) );
  XNOR2_X1 U16284 ( .A(n14489), .B(n14501), .ZN(n14485) );
  OR2_X1 U16285 ( .A1(n14485), .A2(n14924), .ZN(n14625) );
  NOR2_X1 U16286 ( .A1(n14625), .A2(n14486), .ZN(n14487) );
  AOI211_X1 U16287 ( .C1(n14733), .C2(n14489), .A(n14488), .B(n14487), .ZN(
        n14490) );
  OAI211_X1 U16288 ( .C1(n14630), .C2(n14546), .A(n14491), .B(n14490), .ZN(
        P1_U3274) );
  XOR2_X1 U16289 ( .A(n14492), .B(n14495), .Z(n14500) );
  OAI22_X1 U16290 ( .A1(n14494), .A2(n14637), .B1(n14493), .B2(n14517), .ZN(
        n14499) );
  XNOR2_X1 U16291 ( .A(n14496), .B(n14495), .ZN(n14635) );
  NOR2_X1 U16292 ( .A1(n14635), .A2(n14497), .ZN(n14498) );
  AOI211_X1 U16293 ( .C1(n14500), .C2(n14832), .A(n14499), .B(n14498), .ZN(
        n14634) );
  INV_X1 U16294 ( .A(n14501), .ZN(n14502) );
  AOI211_X1 U16295 ( .C1(n14632), .C2(n14520), .A(n14924), .B(n14502), .ZN(
        n14631) );
  INV_X1 U16296 ( .A(n14503), .ZN(n14504) );
  AOI22_X1 U16297 ( .A1(n14743), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14504), 
        .B2(n14732), .ZN(n14505) );
  OAI21_X1 U16298 ( .B1(n14507), .B2(n14506), .A(n14505), .ZN(n14510) );
  NOR2_X1 U16299 ( .A1(n14635), .A2(n14508), .ZN(n14509) );
  AOI211_X1 U16300 ( .C1(n14631), .C2(n14739), .A(n14510), .B(n14509), .ZN(
        n14511) );
  OAI21_X1 U16301 ( .B1(n14634), .B2(n14743), .A(n14511), .ZN(P1_U3275) );
  XOR2_X1 U16302 ( .A(n14514), .B(n14512), .Z(n14644) );
  OAI211_X1 U16303 ( .C1(n14515), .C2(n14514), .A(n14513), .B(n14832), .ZN(
        n14516) );
  OAI21_X1 U16304 ( .B1(n14518), .B2(n14517), .A(n14516), .ZN(n14642) );
  AOI21_X1 U16305 ( .B1(n14519), .B2(n14636), .A(n14924), .ZN(n14521) );
  AND2_X1 U16306 ( .A1(n14521), .A2(n14520), .ZN(n14641) );
  NAND2_X1 U16307 ( .A1(n14641), .A2(n14739), .ZN(n14528) );
  NOR2_X1 U16308 ( .A1(n14522), .A2(n14541), .ZN(n14523) );
  AOI21_X1 U16309 ( .B1(n14743), .B2(P1_REG2_REG_17__SCAN_IN), .A(n14523), 
        .ZN(n14524) );
  OAI21_X1 U16310 ( .B1(n14525), .B2(n14638), .A(n14524), .ZN(n14526) );
  AOI21_X1 U16311 ( .B1(n14636), .B2(n14733), .A(n14526), .ZN(n14527) );
  NAND2_X1 U16312 ( .A1(n14528), .A2(n14527), .ZN(n14529) );
  AOI21_X1 U16313 ( .B1(n14642), .B2(n14544), .A(n14529), .ZN(n14530) );
  OAI21_X1 U16314 ( .B1(n14644), .B2(n14546), .A(n14530), .ZN(P1_U3276) );
  INV_X1 U16315 ( .A(n14531), .ZN(n14533) );
  AOI211_X1 U16316 ( .C1(n14653), .C2(n14533), .A(n14924), .B(n14532), .ZN(
        n14652) );
  XNOR2_X1 U16317 ( .A(n14535), .B(n14534), .ZN(n14538) );
  INV_X1 U16318 ( .A(n14536), .ZN(n14537) );
  AOI21_X1 U16319 ( .B1(n14538), .B2(n14832), .A(n14537), .ZN(n14655) );
  INV_X1 U16320 ( .A(n14655), .ZN(n14539) );
  AOI21_X1 U16321 ( .B1(n14652), .B2(n14540), .A(n14539), .ZN(n14550) );
  INV_X1 U16322 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n14543) );
  OAI22_X1 U16323 ( .A1(n14544), .A2(n14543), .B1(n14542), .B2(n14541), .ZN(
        n14548) );
  XNOR2_X1 U16324 ( .A(n14545), .B(n11181), .ZN(n14656) );
  NOR2_X1 U16325 ( .A1(n14656), .A2(n14546), .ZN(n14547) );
  AOI211_X1 U16326 ( .C1(n14733), .C2(n14653), .A(n14548), .B(n14547), .ZN(
        n14549) );
  OAI21_X1 U16327 ( .B1(n14743), .B2(n14550), .A(n14549), .ZN(P1_U3278) );
  OAI211_X1 U16328 ( .C1(n14552), .C2(n14949), .A(n14551), .B(n14553), .ZN(
        n14657) );
  MUX2_X1 U16329 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14657), .S(n14986), .Z(
        P1_U3559) );
  OAI211_X1 U16330 ( .C1(n14555), .C2(n14949), .A(n14554), .B(n14553), .ZN(
        n14658) );
  MUX2_X1 U16331 ( .A(n14658), .B(P1_REG1_REG_30__SCAN_IN), .S(n14984), .Z(
        P1_U3558) );
  OAI211_X1 U16332 ( .C1(n14559), .C2(n14949), .A(n14558), .B(n14557), .ZN(
        n14560) );
  INV_X1 U16333 ( .A(n14560), .ZN(n14561) );
  AOI22_X1 U16334 ( .A1(n14567), .A2(n14736), .B1(n14566), .B2(n14961), .ZN(
        n14568) );
  OAI211_X1 U16335 ( .C1(n14570), .C2(n14969), .A(n14569), .B(n14568), .ZN(
        n14660) );
  MUX2_X1 U16336 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14660), .S(n14986), .Z(
        P1_U3556) );
  AOI21_X1 U16337 ( .B1(n14572), .B2(n14961), .A(n14571), .ZN(n14573) );
  OAI211_X1 U16338 ( .C1(n14575), .C2(n14966), .A(n14574), .B(n14573), .ZN(
        n14661) );
  MUX2_X1 U16339 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14661), .S(n14986), .Z(
        P1_U3555) );
  AOI211_X1 U16340 ( .C1(n14578), .C2(n14961), .A(n14577), .B(n14576), .ZN(
        n14581) );
  NAND2_X1 U16341 ( .A1(n14579), .A2(n14832), .ZN(n14580) );
  OAI211_X1 U16342 ( .C1(n14969), .C2(n14582), .A(n14581), .B(n14580), .ZN(
        n14662) );
  MUX2_X1 U16343 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14662), .S(n14986), .Z(
        P1_U3554) );
  NAND2_X1 U16344 ( .A1(n14583), .A2(n14927), .ZN(n14588) );
  AOI211_X1 U16345 ( .C1(n14586), .C2(n14961), .A(n14585), .B(n14584), .ZN(
        n14587) );
  OAI211_X1 U16346 ( .C1(n14724), .C2(n14589), .A(n14588), .B(n14587), .ZN(
        n14663) );
  MUX2_X1 U16347 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14663), .S(n14986), .Z(
        P1_U3553) );
  INV_X1 U16348 ( .A(n14966), .ZN(n14945) );
  NAND2_X1 U16349 ( .A1(n14590), .A2(n14945), .ZN(n14593) );
  NAND3_X1 U16350 ( .A1(n14593), .A2(n14592), .A3(n14591), .ZN(n14594) );
  NOR2_X1 U16351 ( .A1(n14595), .A2(n14594), .ZN(n14664) );
  MUX2_X1 U16352 ( .A(n14596), .B(n14664), .S(n14986), .Z(n14597) );
  INV_X1 U16353 ( .A(n14597), .ZN(P1_U3552) );
  NOR4_X1 U16354 ( .A1(n14601), .A2(n14600), .A3(n14599), .A4(n14598), .ZN(
        n14602) );
  OAI21_X1 U16355 ( .B1(n14969), .B2(n14603), .A(n14602), .ZN(n14667) );
  MUX2_X1 U16356 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14667), .S(n14986), .Z(
        P1_U3551) );
  OAI211_X1 U16357 ( .C1(n14949), .C2(n14606), .A(n14605), .B(n14604), .ZN(
        n14607) );
  AOI21_X1 U16358 ( .B1(n14608), .B2(n14927), .A(n14607), .ZN(n14609) );
  OAI21_X1 U16359 ( .B1(n14610), .B2(n14724), .A(n14609), .ZN(n14668) );
  MUX2_X1 U16360 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14668), .S(n14986), .Z(
        P1_U3550) );
  NAND2_X1 U16361 ( .A1(n14611), .A2(n14927), .ZN(n14613) );
  OAI211_X1 U16362 ( .C1(n14614), .C2(n14949), .A(n14613), .B(n14612), .ZN(
        n14615) );
  MUX2_X1 U16363 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14669), .S(n14986), .Z(
        P1_U3549) );
  OAI21_X1 U16364 ( .B1(n14618), .B2(n14949), .A(n14617), .ZN(n14619) );
  AOI211_X1 U16365 ( .C1(n14621), .C2(n14927), .A(n14620), .B(n14619), .ZN(
        n14622) );
  OAI21_X1 U16366 ( .B1(n14724), .B2(n14623), .A(n14622), .ZN(n14670) );
  MUX2_X1 U16367 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14670), .S(n14986), .Z(
        P1_U3548) );
  OAI211_X1 U16368 ( .C1(n14626), .C2(n14949), .A(n14625), .B(n14624), .ZN(
        n14627) );
  AOI21_X1 U16369 ( .B1(n14628), .B2(n14832), .A(n14627), .ZN(n14629) );
  OAI21_X1 U16370 ( .B1(n14969), .B2(n14630), .A(n14629), .ZN(n14671) );
  MUX2_X1 U16371 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14671), .S(n14986), .Z(
        P1_U3547) );
  AOI21_X1 U16372 ( .B1(n14632), .B2(n14961), .A(n14631), .ZN(n14633) );
  OAI211_X1 U16373 ( .C1(n14966), .C2(n14635), .A(n14634), .B(n14633), .ZN(
        n14672) );
  MUX2_X1 U16374 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14672), .S(n14986), .Z(
        P1_U3546) );
  INV_X1 U16375 ( .A(n14636), .ZN(n14639) );
  OAI22_X1 U16376 ( .A1(n14639), .A2(n14949), .B1(n14638), .B2(n14637), .ZN(
        n14640) );
  NOR3_X1 U16377 ( .A1(n14642), .A2(n14641), .A3(n14640), .ZN(n14643) );
  OAI21_X1 U16378 ( .B1(n14969), .B2(n14644), .A(n14643), .ZN(n14673) );
  MUX2_X1 U16379 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14673), .S(n14986), .Z(
        P1_U3545) );
  OAI211_X1 U16380 ( .C1(n14647), .C2(n14949), .A(n14646), .B(n14645), .ZN(
        n14648) );
  AOI21_X1 U16381 ( .B1(n14649), .B2(n14832), .A(n14648), .ZN(n14650) );
  OAI21_X1 U16382 ( .B1(n14651), .B2(n14969), .A(n14650), .ZN(n14674) );
  MUX2_X1 U16383 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14674), .S(n14986), .Z(
        P1_U3544) );
  AOI21_X1 U16384 ( .B1(n14653), .B2(n14961), .A(n14652), .ZN(n14654) );
  OAI211_X1 U16385 ( .C1(n14969), .C2(n14656), .A(n14655), .B(n14654), .ZN(
        n14675) );
  MUX2_X1 U16386 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n14675), .S(n14986), .Z(
        P1_U3543) );
  MUX2_X1 U16387 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14657), .S(n14977), .Z(
        P1_U3527) );
  MUX2_X1 U16388 ( .A(n14658), .B(P1_REG0_REG_30__SCAN_IN), .S(n14975), .Z(
        P1_U3526) );
  MUX2_X1 U16389 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14660), .S(n14977), .Z(
        P1_U3524) );
  MUX2_X1 U16390 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14661), .S(n14977), .Z(
        P1_U3523) );
  MUX2_X1 U16391 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14662), .S(n14977), .Z(
        P1_U3522) );
  MUX2_X1 U16392 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14663), .S(n14977), .Z(
        P1_U3521) );
  MUX2_X1 U16393 ( .A(n14665), .B(n14664), .S(n14977), .Z(n14666) );
  INV_X1 U16394 ( .A(n14666), .ZN(P1_U3520) );
  MUX2_X1 U16395 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14667), .S(n14977), .Z(
        P1_U3519) );
  MUX2_X1 U16396 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14668), .S(n14977), .Z(
        P1_U3518) );
  MUX2_X1 U16397 ( .A(n14669), .B(P1_REG0_REG_21__SCAN_IN), .S(n14975), .Z(
        P1_U3517) );
  MUX2_X1 U16398 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14670), .S(n14977), .Z(
        P1_U3516) );
  MUX2_X1 U16399 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14671), .S(n14977), .Z(
        P1_U3515) );
  MUX2_X1 U16400 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14672), .S(n14953), .Z(
        P1_U3513) );
  MUX2_X1 U16401 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14673), .S(n14953), .Z(
        P1_U3510) );
  MUX2_X1 U16402 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14674), .S(n14953), .Z(
        P1_U3507) );
  MUX2_X1 U16403 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14675), .S(n14953), .Z(
        P1_U3504) );
  NOR4_X1 U16404 ( .A1(n14677), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n14676), .ZN(n14678) );
  AOI21_X1 U16405 ( .B1(n14691), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14678), 
        .ZN(n14679) );
  OAI21_X1 U16406 ( .B1(n14680), .B2(n14694), .A(n14679), .ZN(P1_U3324) );
  INV_X1 U16407 ( .A(n11488), .ZN(n14682) );
  OAI222_X1 U16408 ( .A1(n14683), .A2(P1_U3086), .B1(n14694), .B2(n14682), 
        .C1(n14681), .C2(n14684), .ZN(P1_U3327) );
  OAI222_X1 U16409 ( .A1(P1_U3086), .A2(n6663), .B1(n14694), .B2(n14686), .C1(
        n14685), .C2(n14684), .ZN(P1_U3328) );
  OAI222_X1 U16410 ( .A1(P1_U3086), .A2(n14690), .B1(n14689), .B2(n14688), 
        .C1(n14694), .C2(n14687), .ZN(P1_U3329) );
  AOI22_X1 U16411 ( .A1(n14692), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n14691), .ZN(n14693) );
  OAI21_X1 U16412 ( .B1(n14695), .B2(n14694), .A(n14693), .ZN(P1_U3330) );
  MUX2_X1 U16413 ( .A(n14696), .B(n8784), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16414 ( .A(n14697), .ZN(n14698) );
  MUX2_X1 U16415 ( .A(n14698), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  OAI21_X1 U16416 ( .B1(n14701), .B2(n14700), .A(n14699), .ZN(n14702) );
  XNOR2_X1 U16417 ( .A(n14702), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16418 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14703) );
  OAI21_X1 U16419 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14703), 
        .ZN(U28) );
  AOI21_X1 U16420 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14704) );
  OAI21_X1 U16421 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14704), 
        .ZN(U29) );
  OAI21_X1 U16422 ( .B1(n14707), .B2(n14706), .A(n14705), .ZN(n14708) );
  XNOR2_X1 U16423 ( .A(n14708), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16424 ( .B1(n14711), .B2(n14710), .A(n14709), .ZN(SUB_1596_U57) );
  OAI21_X1 U16425 ( .B1(n14713), .B2(n15044), .A(n14712), .ZN(SUB_1596_U55) );
  AOI21_X1 U16426 ( .B1(n14716), .B2(n14715), .A(n14714), .ZN(SUB_1596_U54) );
  AOI21_X1 U16427 ( .B1(n14719), .B2(n14718), .A(n14717), .ZN(n14720) );
  XOR2_X1 U16428 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14720), .Z(SUB_1596_U70)
         );
  XNOR2_X1 U16429 ( .A(n14721), .B(n14726), .ZN(n14749) );
  INV_X1 U16430 ( .A(n14722), .ZN(n14723) );
  AOI211_X1 U16431 ( .C1(n14726), .C2(n14725), .A(n14724), .B(n14723), .ZN(
        n14727) );
  AOI211_X1 U16432 ( .C1(n14729), .C2(n14749), .A(n14728), .B(n14727), .ZN(
        n14746) );
  INV_X1 U16433 ( .A(n14730), .ZN(n14731) );
  AOI222_X1 U16434 ( .A1(n14734), .A2(n14733), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n14743), .C1(n14732), .C2(n14731), .ZN(n14742) );
  OAI211_X1 U16435 ( .C1(n14745), .C2(n14737), .A(n14736), .B(n14735), .ZN(
        n14744) );
  INV_X1 U16436 ( .A(n14744), .ZN(n14738) );
  AOI22_X1 U16437 ( .A1(n14749), .A2(n14740), .B1(n14739), .B2(n14738), .ZN(
        n14741) );
  OAI211_X1 U16438 ( .C1(n14743), .C2(n14746), .A(n14742), .B(n14741), .ZN(
        P1_U3281) );
  OAI21_X1 U16439 ( .B1(n14745), .B2(n14949), .A(n14744), .ZN(n14748) );
  INV_X1 U16440 ( .A(n14746), .ZN(n14747) );
  AOI211_X1 U16441 ( .C1(n14945), .C2(n14749), .A(n14748), .B(n14747), .ZN(
        n14751) );
  AOI22_X1 U16442 ( .A1(n14953), .A2(n14751), .B1(n10519), .B2(n14975), .ZN(
        P1_U3495) );
  AOI22_X1 U16443 ( .A1(n14986), .A2(n14751), .B1(n14750), .B2(n14984), .ZN(
        P1_U3540) );
  OAI21_X1 U16444 ( .B1(n14754), .B2(n14753), .A(n14752), .ZN(SUB_1596_U63) );
  NOR2_X1 U16445 ( .A1(n14755), .A2(n15226), .ZN(n14784) );
  AOI22_X1 U16446 ( .A1(P3_REG2_REG_13__SCAN_IN), .A2(n15206), .B1(n14770), 
        .B2(n14784), .ZN(n14767) );
  INV_X1 U16447 ( .A(n14779), .ZN(n15162) );
  XNOR2_X1 U16448 ( .A(n14757), .B(n14756), .ZN(n14785) );
  INV_X1 U16449 ( .A(n14785), .ZN(n14764) );
  XNOR2_X1 U16450 ( .A(n13256), .B(n14758), .ZN(n14763) );
  NAND2_X1 U16451 ( .A1(n14759), .A2(n15195), .ZN(n14760) );
  OAI21_X1 U16452 ( .B1(n14775), .B2(n14778), .A(n14760), .ZN(n14761) );
  AOI21_X1 U16453 ( .B1(n14763), .B2(n14762), .A(n14761), .ZN(n14787) );
  OAI21_X1 U16454 ( .B1(n15162), .B2(n14764), .A(n14787), .ZN(n14765) );
  NAND2_X1 U16455 ( .A1(n14765), .A2(n15204), .ZN(n14766) );
  OAI211_X1 U16456 ( .C1(n14768), .C2(n15169), .A(n14767), .B(n14766), .ZN(
        P3_U3220) );
  NOR2_X1 U16457 ( .A1(n14769), .A2(n15226), .ZN(n14796) );
  AOI22_X1 U16458 ( .A1(P3_REG2_REG_11__SCAN_IN), .A2(n15206), .B1(n14770), 
        .B2(n14796), .ZN(n14782) );
  OAI21_X1 U16459 ( .B1(n6550), .B2(n8056), .A(n14771), .ZN(n14797) );
  XNOR2_X1 U16460 ( .A(n14773), .B(n14772), .ZN(n14774) );
  OAI222_X1 U16461 ( .A1(n14778), .A2(n14777), .B1(n14776), .B2(n14775), .C1(
        n14774), .C2(n15198), .ZN(n14795) );
  AOI21_X1 U16462 ( .B1(n14779), .B2(n14797), .A(n14795), .ZN(n14780) );
  OR2_X1 U16463 ( .A1(n14780), .A2(n15206), .ZN(n14781) );
  OAI211_X1 U16464 ( .C1(n14783), .C2(n15169), .A(n14782), .B(n14781), .ZN(
        P3_U3222) );
  AOI21_X1 U16465 ( .B1(n14785), .B2(n14798), .A(n14784), .ZN(n14786) );
  INV_X1 U16466 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14788) );
  AOI22_X1 U16467 ( .A1(n15240), .A2(n14800), .B1(n14788), .B2(n15241), .ZN(
        P3_U3472) );
  OAI22_X1 U16468 ( .A1(n14791), .A2(n14790), .B1(n14789), .B2(n15226), .ZN(
        n14792) );
  NOR2_X1 U16469 ( .A1(n14793), .A2(n14792), .ZN(n14802) );
  AOI22_X1 U16470 ( .A1(n15240), .A2(n14802), .B1(n14794), .B2(n15241), .ZN(
        P3_U3471) );
  AOI211_X1 U16471 ( .C1(n14798), .C2(n14797), .A(n14796), .B(n14795), .ZN(
        n14804) );
  INV_X1 U16472 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14799) );
  AOI22_X1 U16473 ( .A1(n15240), .A2(n14804), .B1(n14799), .B2(n15241), .ZN(
        P3_U3470) );
  INV_X1 U16474 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14801) );
  AOI22_X1 U16475 ( .A1(n15234), .A2(n14801), .B1(n14800), .B2(n15232), .ZN(
        P3_U3429) );
  INV_X1 U16476 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14803) );
  AOI22_X1 U16477 ( .A1(n15234), .A2(n14803), .B1(n14802), .B2(n15232), .ZN(
        P3_U3426) );
  INV_X1 U16478 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14805) );
  AOI22_X1 U16479 ( .A1(n15234), .A2(n14805), .B1(n14804), .B2(n15232), .ZN(
        P3_U3423) );
  AND2_X1 U16480 ( .A1(n14806), .A2(n14961), .ZN(n14972) );
  OAI22_X1 U16481 ( .A1(n14808), .A2(n14871), .B1(n14870), .B2(n14807), .ZN(
        n14814) );
  OAI211_X1 U16482 ( .C1(n14811), .C2(n14810), .A(n14822), .B(n14809), .ZN(
        n14812) );
  INV_X1 U16483 ( .A(n14812), .ZN(n14813) );
  AOI211_X1 U16484 ( .C1(n14972), .C2(n14815), .A(n14814), .B(n14813), .ZN(
        n14817) );
  OAI211_X1 U16485 ( .C1(n14883), .C2(n14818), .A(n14817), .B(n14816), .ZN(
        P1_U3217) );
  OAI22_X1 U16486 ( .A1(n14819), .A2(n14871), .B1(n14870), .B2(n14872), .ZN(
        n14827) );
  AOI21_X1 U16487 ( .B1(n14822), .B2(n14821), .A(n14820), .ZN(n14823) );
  INV_X1 U16488 ( .A(n14823), .ZN(n14825) );
  AOI21_X1 U16489 ( .B1(n14825), .B2(n14824), .A(n14875), .ZN(n14826) );
  AOI211_X1 U16490 ( .C1(n14879), .C2(n14828), .A(n14827), .B(n14826), .ZN(
        n14830) );
  OAI211_X1 U16491 ( .C1(n14883), .C2(n14831), .A(n14830), .B(n14829), .ZN(
        P1_U3236) );
  NAND3_X1 U16492 ( .A1(n14833), .A2(n14832), .A3(n10974), .ZN(n14838) );
  AOI21_X1 U16493 ( .B1(n14835), .B2(n14961), .A(n14834), .ZN(n14837) );
  NAND3_X1 U16494 ( .A1(n14838), .A2(n14837), .A3(n14836), .ZN(n14839) );
  AOI21_X1 U16495 ( .B1(n14840), .B2(n14927), .A(n14839), .ZN(n14842) );
  AOI22_X1 U16496 ( .A1(n14986), .A2(n14842), .B1(n10843), .B2(n14984), .ZN(
        P1_U3541) );
  INV_X1 U16497 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14841) );
  AOI22_X1 U16498 ( .A1(n14953), .A2(n14842), .B1(n14841), .B2(n14975), .ZN(
        P1_U3498) );
  OAI21_X1 U16499 ( .B1(n14845), .B2(n14844), .A(n14843), .ZN(n14846) );
  XNOR2_X1 U16500 ( .A(n14846), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  AOI21_X1 U16501 ( .B1(n14849), .B2(n14848), .A(n14847), .ZN(n14850) );
  XOR2_X1 U16502 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n14850), .Z(SUB_1596_U68)
         );
  AOI21_X1 U16503 ( .B1(n14853), .B2(n14852), .A(n14851), .ZN(n14854) );
  XOR2_X1 U16504 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n14854), .Z(SUB_1596_U67)
         );
  OAI222_X1 U16505 ( .A1(n14859), .A2(n14858), .B1(n14859), .B2(n14857), .C1(
        n14856), .C2(n14855), .ZN(SUB_1596_U66) );
  OAI222_X1 U16506 ( .A1(n14864), .A2(n14863), .B1(n14864), .B2(n14862), .C1(
        n14861), .C2(n14860), .ZN(SUB_1596_U65) );
  AOI21_X1 U16507 ( .B1(n14867), .B2(n14866), .A(n14865), .ZN(n14868) );
  XOR2_X1 U16508 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14868), .Z(SUB_1596_U64)
         );
  OAI22_X1 U16509 ( .A1(n14872), .A2(n14871), .B1(n14870), .B2(n14869), .ZN(
        n14878) );
  XOR2_X1 U16510 ( .A(n14873), .B(n14874), .Z(n14876) );
  NOR2_X1 U16511 ( .A1(n14876), .A2(n14875), .ZN(n14877) );
  AOI211_X1 U16512 ( .C1(n14879), .C2(n14962), .A(n14878), .B(n14877), .ZN(
        n14881) );
  OAI211_X1 U16513 ( .C1(n14883), .C2(n14882), .A(n14881), .B(n14880), .ZN(
        P1_U3231) );
  AND2_X1 U16514 ( .A1(n6663), .A2(n14884), .ZN(n14888) );
  NOR2_X1 U16515 ( .A1(n14886), .A2(n14888), .ZN(n14887) );
  MUX2_X1 U16516 ( .A(n14888), .B(n14887), .S(P1_IR_REG_0__SCAN_IN), .Z(n14890) );
  OR2_X1 U16517 ( .A1(n14890), .A2(n14889), .ZN(n14893) );
  AOI22_X1 U16518 ( .A1(n14891), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14892) );
  OAI21_X1 U16519 ( .B1(n14894), .B2(n14893), .A(n14892), .ZN(P1_U3243) );
  AOI21_X1 U16520 ( .B1(n14896), .B2(P1_REG2_REG_15__SCAN_IN), .A(n14895), 
        .ZN(n14907) );
  OAI21_X1 U16521 ( .B1(n14899), .B2(n14898), .A(n14897), .ZN(n14900) );
  NAND2_X1 U16522 ( .A1(n14901), .A2(n14900), .ZN(n14905) );
  NAND2_X1 U16523 ( .A1(n14903), .A2(n14902), .ZN(n14904) );
  OAI211_X1 U16524 ( .C1(n14907), .C2(n14906), .A(n14905), .B(n14904), .ZN(
        n14908) );
  INV_X1 U16525 ( .A(n14908), .ZN(n14910) );
  OAI211_X1 U16526 ( .C1(n14912), .C2(n14911), .A(n14910), .B(n14909), .ZN(
        P1_U3258) );
  AND2_X1 U16527 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14917), .ZN(P1_U3294) );
  AND2_X1 U16528 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14917), .ZN(P1_U3295) );
  AND2_X1 U16529 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14917), .ZN(P1_U3296) );
  AND2_X1 U16530 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14917), .ZN(P1_U3297) );
  INV_X1 U16531 ( .A(n14917), .ZN(n14916) );
  NOR2_X1 U16532 ( .A1(n14916), .A2(n14913), .ZN(P1_U3298) );
  AND2_X1 U16533 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14917), .ZN(P1_U3299) );
  AND2_X1 U16534 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14917), .ZN(P1_U3300) );
  AND2_X1 U16535 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14917), .ZN(P1_U3301) );
  AND2_X1 U16536 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14917), .ZN(P1_U3302) );
  AND2_X1 U16537 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14917), .ZN(P1_U3303) );
  AND2_X1 U16538 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14917), .ZN(P1_U3304) );
  AND2_X1 U16539 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14917), .ZN(P1_U3305) );
  NOR2_X1 U16540 ( .A1(n14916), .A2(n14914), .ZN(P1_U3306) );
  AND2_X1 U16541 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14917), .ZN(P1_U3307) );
  AND2_X1 U16542 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14917), .ZN(P1_U3308) );
  AND2_X1 U16543 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14917), .ZN(P1_U3309) );
  AND2_X1 U16544 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14917), .ZN(P1_U3310) );
  AND2_X1 U16545 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14917), .ZN(P1_U3311) );
  AND2_X1 U16546 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14917), .ZN(P1_U3312) );
  AND2_X1 U16547 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14917), .ZN(P1_U3313) );
  AND2_X1 U16548 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14917), .ZN(P1_U3314) );
  AND2_X1 U16549 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14917), .ZN(P1_U3315) );
  AND2_X1 U16550 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14917), .ZN(P1_U3316) );
  AND2_X1 U16551 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14917), .ZN(P1_U3317) );
  AND2_X1 U16552 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14917), .ZN(P1_U3318) );
  AND2_X1 U16553 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14917), .ZN(P1_U3319) );
  AND2_X1 U16554 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14917), .ZN(P1_U3320) );
  AND2_X1 U16555 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14917), .ZN(P1_U3321) );
  NOR2_X1 U16556 ( .A1(n14916), .A2(n14915), .ZN(P1_U3322) );
  AND2_X1 U16557 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14917), .ZN(P1_U3323) );
  AOI22_X1 U16558 ( .A1(n14977), .A2(n14918), .B1(n8694), .B2(n14975), .ZN(
        P1_U3459) );
  INV_X1 U16559 ( .A(n14919), .ZN(n14928) );
  AOI22_X1 U16560 ( .A1(n9387), .A2(n14921), .B1(n14920), .B2(n14961), .ZN(
        n14922) );
  OAI211_X1 U16561 ( .C1(n14925), .C2(n14924), .A(n14923), .B(n14922), .ZN(
        n14926) );
  AOI21_X1 U16562 ( .B1(n14928), .B2(n14927), .A(n14926), .ZN(n14978) );
  INV_X1 U16563 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14929) );
  AOI22_X1 U16564 ( .A1(n14977), .A2(n14978), .B1(n14929), .B2(n14975), .ZN(
        P1_U3462) );
  NAND2_X1 U16565 ( .A1(n14930), .A2(n14945), .ZN(n14932) );
  OAI211_X1 U16566 ( .C1(n14933), .C2(n14949), .A(n14932), .B(n14931), .ZN(
        n14935) );
  NOR2_X1 U16567 ( .A1(n14935), .A2(n14934), .ZN(n14979) );
  INV_X1 U16568 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14936) );
  AOI22_X1 U16569 ( .A1(n14977), .A2(n14979), .B1(n14936), .B2(n14975), .ZN(
        P1_U3465) );
  OAI21_X1 U16570 ( .B1(n14938), .B2(n14949), .A(n14937), .ZN(n14941) );
  INV_X1 U16571 ( .A(n14939), .ZN(n14940) );
  AOI211_X1 U16572 ( .C1(n14945), .C2(n14942), .A(n14941), .B(n14940), .ZN(
        n14980) );
  INV_X1 U16573 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14943) );
  AOI22_X1 U16574 ( .A1(n14953), .A2(n14980), .B1(n14943), .B2(n14975), .ZN(
        P1_U3468) );
  INV_X1 U16575 ( .A(n14944), .ZN(n14950) );
  NAND2_X1 U16576 ( .A1(n14946), .A2(n14945), .ZN(n14948) );
  OAI211_X1 U16577 ( .C1(n14950), .C2(n14949), .A(n14948), .B(n14947), .ZN(
        n14952) );
  NOR2_X1 U16578 ( .A1(n14952), .A2(n14951), .ZN(n14981) );
  AOI22_X1 U16579 ( .A1(n14953), .A2(n14981), .B1(n9312), .B2(n14975), .ZN(
        P1_U3477) );
  AOI211_X1 U16580 ( .C1(n14956), .C2(n14961), .A(n14955), .B(n14954), .ZN(
        n14957) );
  OAI21_X1 U16581 ( .B1(n14969), .B2(n14958), .A(n14957), .ZN(n14959) );
  INV_X1 U16582 ( .A(n14959), .ZN(n14982) );
  AOI22_X1 U16583 ( .A1(n14977), .A2(n14982), .B1(n9930), .B2(n14975), .ZN(
        P1_U3483) );
  AOI21_X1 U16584 ( .B1(n14962), .B2(n14961), .A(n14960), .ZN(n14963) );
  OAI211_X1 U16585 ( .C1(n14966), .C2(n14965), .A(n14964), .B(n14963), .ZN(
        n14967) );
  INV_X1 U16586 ( .A(n14967), .ZN(n14983) );
  INV_X1 U16587 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14968) );
  AOI22_X1 U16588 ( .A1(n14977), .A2(n14983), .B1(n14968), .B2(n14975), .ZN(
        P1_U3486) );
  NOR2_X1 U16589 ( .A1(n14970), .A2(n14969), .ZN(n14974) );
  NOR4_X1 U16590 ( .A1(n14974), .A2(n14973), .A3(n14972), .A4(n14971), .ZN(
        n14985) );
  INV_X1 U16591 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14976) );
  AOI22_X1 U16592 ( .A1(n14977), .A2(n14985), .B1(n14976), .B2(n14975), .ZN(
        P1_U3489) );
  AOI22_X1 U16593 ( .A1(n14986), .A2(n14978), .B1(n8788), .B2(n14984), .ZN(
        P1_U3529) );
  AOI22_X1 U16594 ( .A1(n14986), .A2(n14979), .B1(n8986), .B2(n14984), .ZN(
        P1_U3530) );
  AOI22_X1 U16595 ( .A1(n14986), .A2(n14980), .B1(n8997), .B2(n14984), .ZN(
        P1_U3531) );
  AOI22_X1 U16596 ( .A1(n14986), .A2(n14981), .B1(n9314), .B2(n14984), .ZN(
        P1_U3534) );
  AOI22_X1 U16597 ( .A1(n14986), .A2(n14982), .B1(n9933), .B2(n14984), .ZN(
        P1_U3536) );
  AOI22_X1 U16598 ( .A1(n14986), .A2(n14983), .B1(n10119), .B2(n14984), .ZN(
        P1_U3537) );
  AOI22_X1 U16599 ( .A1(n14986), .A2(n14985), .B1(n10386), .B2(n14984), .ZN(
        P1_U3538) );
  NOR2_X1 U16600 ( .A1(n14987), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16601 ( .A1(n14987), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n15000) );
  OAI21_X1 U16602 ( .B1(n14990), .B2(n14989), .A(n14988), .ZN(n14991) );
  OAI22_X1 U16603 ( .A1(n14993), .A2(n14992), .B1(n15046), .B2(n14991), .ZN(
        n14994) );
  INV_X1 U16604 ( .A(n14994), .ZN(n14999) );
  OAI211_X1 U16605 ( .C1(n14997), .C2(n14996), .A(n15039), .B(n14995), .ZN(
        n14998) );
  NAND3_X1 U16606 ( .A1(n15000), .A2(n14999), .A3(n14998), .ZN(P2_U3216) );
  INV_X1 U16607 ( .A(n15001), .ZN(n15008) );
  OAI211_X1 U16608 ( .C1(n15005), .C2(n15004), .A(n15003), .B(n15002), .ZN(
        n15006) );
  INV_X1 U16609 ( .A(n15006), .ZN(n15007) );
  AOI211_X1 U16610 ( .C1(n15052), .C2(n15009), .A(n15008), .B(n15007), .ZN(
        n15014) );
  OAI211_X1 U16611 ( .C1(n15012), .C2(n15011), .A(n15039), .B(n15010), .ZN(
        n15013) );
  OAI211_X1 U16612 ( .C1(n15061), .C2(n15015), .A(n15014), .B(n15013), .ZN(
        P2_U3218) );
  OAI21_X1 U16613 ( .B1(n15018), .B2(n15017), .A(n15016), .ZN(n15019) );
  OR2_X1 U16614 ( .A1(n15046), .A2(n15019), .ZN(n15021) );
  OAI211_X1 U16615 ( .C1(n15034), .C2(n15022), .A(n15021), .B(n15020), .ZN(
        n15023) );
  INV_X1 U16616 ( .A(n15023), .ZN(n15028) );
  OAI211_X1 U16617 ( .C1(n15026), .C2(n15025), .A(n15039), .B(n15024), .ZN(
        n15027) );
  OAI211_X1 U16618 ( .C1(n15061), .C2(n15247), .A(n15028), .B(n15027), .ZN(
        P2_U3219) );
  AOI211_X1 U16619 ( .C1(n15031), .C2(n15030), .A(n15046), .B(n15029), .ZN(
        n15036) );
  OAI21_X1 U16620 ( .B1(n15034), .B2(n15033), .A(n15032), .ZN(n15035) );
  NOR2_X1 U16621 ( .A1(n15036), .A2(n15035), .ZN(n15043) );
  INV_X1 U16622 ( .A(n15037), .ZN(n15038) );
  OAI211_X1 U16623 ( .C1(n15041), .C2(n15040), .A(n15039), .B(n15038), .ZN(
        n15042) );
  OAI211_X1 U16624 ( .C1(n15061), .C2(n15044), .A(n15043), .B(n15042), .ZN(
        P2_U3222) );
  INV_X1 U16625 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15060) );
  NOR2_X1 U16626 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10426), .ZN(n15050) );
  AOI211_X1 U16627 ( .C1(n15048), .C2(n15047), .A(n15046), .B(n15045), .ZN(
        n15049) );
  AOI211_X1 U16628 ( .C1(n15052), .C2(n15051), .A(n15050), .B(n15049), .ZN(
        n15059) );
  AOI211_X1 U16629 ( .C1(n15056), .C2(n15055), .A(n15054), .B(n15053), .ZN(
        n15057) );
  INV_X1 U16630 ( .A(n15057), .ZN(n15058) );
  OAI211_X1 U16631 ( .C1(n15061), .C2(n15060), .A(n15059), .B(n15058), .ZN(
        P2_U3227) );
  AOI22_X1 U16632 ( .A1(n15075), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n15063), 
        .B2(n15062), .ZN(n15067) );
  NAND2_X1 U16633 ( .A1(n15065), .A2(n15064), .ZN(n15066) );
  OAI211_X1 U16634 ( .C1(n15069), .C2(n15068), .A(n15067), .B(n15066), .ZN(
        n15070) );
  AOI21_X1 U16635 ( .B1(n15072), .B2(n15071), .A(n15070), .ZN(n15073) );
  OAI21_X1 U16636 ( .B1(n15075), .B2(n15074), .A(n15073), .ZN(P2_U3258) );
  INV_X1 U16637 ( .A(n15087), .ZN(n15082) );
  AND2_X1 U16638 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15081), .ZN(P2_U3266) );
  AND2_X1 U16639 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15081), .ZN(P2_U3267) );
  AND2_X1 U16640 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15081), .ZN(P2_U3268) );
  AND2_X1 U16641 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15081), .ZN(P2_U3269) );
  AND2_X1 U16642 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15081), .ZN(P2_U3270) );
  AND2_X1 U16643 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15081), .ZN(P2_U3271) );
  AND2_X1 U16644 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15081), .ZN(P2_U3272) );
  AND2_X1 U16645 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15081), .ZN(P2_U3273) );
  NOR2_X1 U16646 ( .A1(n15080), .A2(n15077), .ZN(P2_U3274) );
  AND2_X1 U16647 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15081), .ZN(P2_U3275) );
  AND2_X1 U16648 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15081), .ZN(P2_U3276) );
  AND2_X1 U16649 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15081), .ZN(P2_U3277) );
  AND2_X1 U16650 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15081), .ZN(P2_U3278) );
  AND2_X1 U16651 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15081), .ZN(P2_U3279) );
  AND2_X1 U16652 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15081), .ZN(P2_U3280) );
  AND2_X1 U16653 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15081), .ZN(P2_U3281) );
  AND2_X1 U16654 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15081), .ZN(P2_U3282) );
  AND2_X1 U16655 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15081), .ZN(P2_U3283) );
  AND2_X1 U16656 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15081), .ZN(P2_U3284) );
  NOR2_X1 U16657 ( .A1(n15080), .A2(n15078), .ZN(P2_U3285) );
  AND2_X1 U16658 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15081), .ZN(P2_U3286) );
  NOR2_X1 U16659 ( .A1(n15080), .A2(n15079), .ZN(P2_U3287) );
  AND2_X1 U16660 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15081), .ZN(P2_U3288) );
  AND2_X1 U16661 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15081), .ZN(P2_U3289) );
  AND2_X1 U16662 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15081), .ZN(P2_U3290) );
  AND2_X1 U16663 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15081), .ZN(P2_U3291) );
  AND2_X1 U16664 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15081), .ZN(P2_U3292) );
  AND2_X1 U16665 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15081), .ZN(P2_U3293) );
  AND2_X1 U16666 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15081), .ZN(P2_U3294) );
  AND2_X1 U16667 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15081), .ZN(P2_U3295) );
  AOI22_X1 U16668 ( .A1(n15087), .A2(n15084), .B1(n15083), .B2(n15082), .ZN(
        P2_U3416) );
  OAI21_X1 U16669 ( .B1(n15087), .B2(n15086), .A(n15085), .ZN(P2_U3417) );
  AOI21_X1 U16670 ( .B1(n15098), .B2(n15089), .A(n15088), .ZN(n15091) );
  OAI211_X1 U16671 ( .C1(n15093), .C2(n15092), .A(n15091), .B(n15090), .ZN(
        n15094) );
  INV_X1 U16672 ( .A(n15094), .ZN(n15108) );
  INV_X1 U16673 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15095) );
  AOI22_X1 U16674 ( .A1(n15106), .A2(n15108), .B1(n15095), .B2(n15104), .ZN(
        P2_U3442) );
  AOI21_X1 U16675 ( .B1(n15098), .B2(n15097), .A(n15096), .ZN(n15099) );
  OAI211_X1 U16676 ( .C1(n15102), .C2(n15101), .A(n15100), .B(n15099), .ZN(
        n15103) );
  INV_X1 U16677 ( .A(n15103), .ZN(n15111) );
  INV_X1 U16678 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15105) );
  AOI22_X1 U16679 ( .A1(n15106), .A2(n15111), .B1(n15105), .B2(n15104), .ZN(
        P2_U3448) );
  AOI22_X1 U16680 ( .A1(n15112), .A2(n15108), .B1(n15107), .B2(n15109), .ZN(
        P2_U3503) );
  AOI22_X1 U16681 ( .A1(n15112), .A2(n15111), .B1(n15110), .B2(n15109), .ZN(
        P2_U3505) );
  NOR2_X1 U16682 ( .A1(P3_U3897), .A2(n15113), .ZN(P3_U3150) );
  MUX2_X1 U16683 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n9963), .S(n15127), .Z(
        n15116) );
  NAND2_X1 U16684 ( .A1(n15115), .A2(n15116), .ZN(n15114) );
  OAI21_X1 U16685 ( .B1(n15116), .B2(n15115), .A(n15114), .ZN(n15130) );
  AOI21_X1 U16686 ( .B1(n15119), .B2(n15118), .A(n15117), .ZN(n15120) );
  NOR2_X1 U16687 ( .A1(n15140), .A2(n15120), .ZN(n15129) );
  AND3_X1 U16688 ( .A1(n15123), .A2(n15122), .A3(n15121), .ZN(n15124) );
  OAI21_X1 U16689 ( .B1(n15125), .B2(n15124), .A(n15146), .ZN(n15126) );
  OAI21_X1 U16690 ( .B1(n15150), .B2(n15127), .A(n15126), .ZN(n15128) );
  AOI211_X1 U16691 ( .C1(n15154), .C2(n15130), .A(n15129), .B(n15128), .ZN(
        n15132) );
  OAI211_X1 U16692 ( .C1(n15133), .C2(n15157), .A(n15132), .B(n15131), .ZN(
        P3_U3188) );
  INV_X1 U16693 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15158) );
  MUX2_X1 U16694 ( .A(P3_REG2_REG_8__SCAN_IN), .B(n10161), .S(n15149), .Z(
        n15136) );
  NAND2_X1 U16695 ( .A1(n15135), .A2(n15136), .ZN(n15134) );
  OAI21_X1 U16696 ( .B1(n15136), .B2(n15135), .A(n15134), .ZN(n15153) );
  INV_X1 U16697 ( .A(n15137), .ZN(n15139) );
  NAND2_X1 U16698 ( .A1(n15139), .A2(n15138), .ZN(n15142) );
  AOI21_X1 U16699 ( .B1(n15142), .B2(n15141), .A(n15140), .ZN(n15152) );
  OAI21_X1 U16700 ( .B1(n15145), .B2(n15144), .A(n15143), .ZN(n15147) );
  NAND2_X1 U16701 ( .A1(n15147), .A2(n15146), .ZN(n15148) );
  OAI21_X1 U16702 ( .B1(n15150), .B2(n15149), .A(n15148), .ZN(n15151) );
  AOI211_X1 U16703 ( .C1(n15154), .C2(n15153), .A(n15152), .B(n15151), .ZN(
        n15156) );
  OAI211_X1 U16704 ( .C1(n15158), .C2(n15157), .A(n15156), .B(n15155), .ZN(
        P3_U3190) );
  INV_X1 U16705 ( .A(n15159), .ZN(n15161) );
  OAI21_X1 U16706 ( .B1(n15162), .B2(n15161), .A(n15160), .ZN(n15167) );
  INV_X1 U16707 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15163) );
  OAI22_X1 U16708 ( .A1(n15165), .A2(n15164), .B1(n15163), .B2(n15204), .ZN(
        n15166) );
  AOI21_X1 U16709 ( .B1(n15167), .B2(n15204), .A(n15166), .ZN(n15168) );
  OAI21_X1 U16710 ( .B1(n15170), .B2(n15169), .A(n15168), .ZN(P3_U3224) );
  XNOR2_X1 U16711 ( .A(n15171), .B(n15175), .ZN(n15180) );
  AOI22_X1 U16712 ( .A1(n15173), .A2(n15192), .B1(n15195), .B2(n15172), .ZN(
        n15179) );
  OAI21_X1 U16713 ( .B1(n15176), .B2(n15175), .A(n15174), .ZN(n15213) );
  INV_X1 U16714 ( .A(n15177), .ZN(n15191) );
  NAND2_X1 U16715 ( .A1(n15213), .A2(n15191), .ZN(n15178) );
  OAI211_X1 U16716 ( .C1(n15180), .C2(n15198), .A(n15179), .B(n15178), .ZN(
        n15211) );
  INV_X1 U16717 ( .A(n15213), .ZN(n15184) );
  NOR2_X1 U16718 ( .A1(n7722), .A2(n15226), .ZN(n15212) );
  INV_X1 U16719 ( .A(n15212), .ZN(n15181) );
  OAI22_X1 U16720 ( .A1(n15184), .A2(n15183), .B1(n15182), .B2(n15181), .ZN(
        n15185) );
  AOI211_X1 U16721 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15201), .A(n15211), .B(
        n15185), .ZN(n15186) );
  AOI22_X1 U16722 ( .A1(n15206), .A2(n9171), .B1(n15186), .B2(n15204), .ZN(
        P3_U3231) );
  NOR2_X1 U16723 ( .A1(n15187), .A2(n15226), .ZN(n15208) );
  XNOR2_X1 U16724 ( .A(n15189), .B(n15188), .ZN(n15199) );
  XNOR2_X1 U16725 ( .A(n15190), .B(n15189), .ZN(n15209) );
  NAND2_X1 U16726 ( .A1(n15209), .A2(n15191), .ZN(n15197) );
  AOI22_X1 U16727 ( .A1(n15195), .A2(n15194), .B1(n15193), .B2(n15192), .ZN(
        n15196) );
  OAI211_X1 U16728 ( .C1(n15199), .C2(n15198), .A(n15197), .B(n15196), .ZN(
        n15207) );
  AOI21_X1 U16729 ( .B1(n15208), .B2(n15200), .A(n15207), .ZN(n15205) );
  AOI22_X1 U16730 ( .A1(n15202), .A2(n15209), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15201), .ZN(n15203) );
  OAI221_X1 U16731 ( .B1(n15206), .B2(n15205), .C1(n15204), .C2(n9174), .A(
        n15203), .ZN(P3_U3232) );
  INV_X1 U16732 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15210) );
  AOI211_X1 U16733 ( .C1(n15223), .C2(n15209), .A(n15208), .B(n15207), .ZN(
        n15235) );
  AOI22_X1 U16734 ( .A1(n15234), .A2(n15210), .B1(n15235), .B2(n15232), .ZN(
        P3_U3393) );
  INV_X1 U16735 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15214) );
  AOI211_X1 U16736 ( .C1(n15223), .C2(n15213), .A(n15212), .B(n15211), .ZN(
        n15236) );
  AOI22_X1 U16737 ( .A1(n15234), .A2(n15214), .B1(n15236), .B2(n15232), .ZN(
        P3_U3396) );
  INV_X1 U16738 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15219) );
  INV_X1 U16739 ( .A(n15215), .ZN(n15218) );
  AOI211_X1 U16740 ( .C1(n15218), .C2(n15223), .A(n15217), .B(n15216), .ZN(
        n15237) );
  AOI22_X1 U16741 ( .A1(n15234), .A2(n15219), .B1(n15237), .B2(n15232), .ZN(
        P3_U3405) );
  INV_X1 U16742 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15225) );
  INV_X1 U16743 ( .A(n15220), .ZN(n15224) );
  AOI211_X1 U16744 ( .C1(n15224), .C2(n15223), .A(n15222), .B(n15221), .ZN(
        n15239) );
  AOI22_X1 U16745 ( .A1(n15234), .A2(n15225), .B1(n15239), .B2(n15232), .ZN(
        P3_U3414) );
  INV_X1 U16746 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15233) );
  OAI22_X1 U16747 ( .A1(n15229), .A2(n15228), .B1(n15227), .B2(n15226), .ZN(
        n15230) );
  NOR2_X1 U16748 ( .A1(n15231), .A2(n15230), .ZN(n15242) );
  AOI22_X1 U16749 ( .A1(n15234), .A2(n15233), .B1(n15242), .B2(n15232), .ZN(
        P3_U3420) );
  AOI22_X1 U16750 ( .A1(n15240), .A2(n15235), .B1(n9161), .B2(n15241), .ZN(
        P3_U3460) );
  AOI22_X1 U16751 ( .A1(n15240), .A2(n15236), .B1(n9158), .B2(n15241), .ZN(
        P3_U3461) );
  AOI22_X1 U16752 ( .A1(n15240), .A2(n15237), .B1(n9374), .B2(n15241), .ZN(
        P3_U3464) );
  AOI22_X1 U16753 ( .A1(n15240), .A2(n15239), .B1(n15238), .B2(n15241), .ZN(
        P3_U3467) );
  AOI22_X1 U16754 ( .A1(n15240), .A2(n15242), .B1(n10347), .B2(n15241), .ZN(
        P3_U3469) );
  AOI21_X1 U16755 ( .B1(n15245), .B2(n15244), .A(n15243), .ZN(SUB_1596_U59) );
  OAI21_X1 U16756 ( .B1(n15248), .B2(n15247), .A(n15246), .ZN(SUB_1596_U58) );
  XOR2_X1 U16757 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15249), .Z(SUB_1596_U53) );
  AOI21_X1 U16758 ( .B1(n15252), .B2(n15251), .A(n15250), .ZN(SUB_1596_U56) );
  AOI21_X1 U16759 ( .B1(n15255), .B2(n15254), .A(n15253), .ZN(n15256) );
  XOR2_X1 U16760 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15256), .Z(SUB_1596_U60) );
  AOI21_X1 U16761 ( .B1(n15259), .B2(n15258), .A(n15257), .ZN(SUB_1596_U5) );
  CLKBUF_X2 U11338 ( .A(n8843), .Z(n12400) );
  NAND2_X2 U7295 ( .A1(n10313), .A2(n12444), .ZN(n13459) );
  AND2_X1 U7305 ( .A1(n11473), .A2(n8602), .ZN(n12489) );
  XNOR2_X1 U7340 ( .A(n11063), .B(n11064), .ZN(n10719) );
  CLKBUF_X1 U8586 ( .A(n12294), .Z(n6593) );
  CLKBUF_X1 U8843 ( .A(n12281), .Z(n6604) );
  CLKBUF_X1 U9314 ( .A(n12110), .Z(n6699) );
  AOI211_X1 U9461 ( .C1(n10060), .C2(n10059), .A(n12739), .B(n6553), .ZN(
        n10061) );
  NAND2_X2 U9505 ( .A1(n9658), .A2(n9657), .ZN(n12739) );
endmodule

