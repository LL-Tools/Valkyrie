

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput63, keyinput62, keyinput61, 
        keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, 
        keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, 
        keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, 
        keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, 
        keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, 
        keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, 
        keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, 
        keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, 
        keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, 
        keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, 
        keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2945, n2946, n2948, n2949, n2951, n2952, n2953, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667;

  AND2_X1 U3393 ( .A1(n5284), .A2(n5283), .ZN(n5285) );
  AND2_X1 U3394 ( .A1(n5452), .A2(n3751), .ZN(n5502) );
  NOR2_X1 U3395 ( .A1(n5492), .A2(n3104), .ZN(n5361) );
  NAND2_X1 U3396 ( .A1(n3306), .A2(n3307), .ZN(n4220) );
  NOR2_X1 U3397 ( .A1(n4691), .A2(n4065), .ZN(n4000) );
  AND2_X2 U3398 ( .A1(n5400), .A2(n2963), .ZN(n3126) );
  CLKBUF_X2 U3399 ( .A(n3313), .Z(n3909) );
  AND2_X1 U3400 ( .A1(n2961), .A2(n5391), .ZN(n3311) );
  BUF_X2 U3401 ( .A(n3179), .Z(n3732) );
  CLKBUF_X2 U3402 ( .A(n3162), .Z(n3823) );
  AND2_X1 U3403 ( .A1(n2959), .A2(n5152), .ZN(n3312) );
  AND2_X1 U3404 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4219) );
  NAND2_X2 U3407 ( .A1(n4288), .A2(n4465), .ZN(n3100) );
  OR2_X1 U3408 ( .A1(n5549), .A2(n5183), .ZN(n5353) );
  INV_X1 U3409 ( .A(n5581), .ZN(n4811) );
  INV_X1 U3410 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6369) );
  XNOR2_X1 U3411 ( .A(n4220), .B(n6309), .ZN(n4523) );
  AND2_X1 U3412 ( .A1(n3327), .A2(n3328), .ZN(n3376) );
  INV_X1 U3413 ( .A(n4121), .ZN(n4092) );
  NOR2_X1 U3414 ( .A1(n4140), .A2(n4152), .ZN(n3458) );
  INV_X1 U3415 ( .A(n5581), .ZN(n5875) );
  NAND2_X1 U3416 ( .A1(n5581), .A2(n4699), .ZN(n4805) );
  NAND2_X1 U3417 ( .A1(n3295), .A2(n3329), .ZN(n4654) );
  NAND2_X1 U3418 ( .A1(n4026), .A2(n4284), .ZN(n4243) );
  INV_X2 U3419 ( .A(n4047), .ZN(n4284) );
  OAI22_X1 U3420 ( .A1(n5337), .A2(n5336), .B1(n5335), .B2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5338) );
  INV_X1 U3421 ( .A(n5958), .ZN(n5997) );
  MUX2_X2 U3422 ( .A(n3395), .B(n3394), .S(n3393), .Z(n4615) );
  OAI21_X1 U3423 ( .B1(n4654), .B2(STATE2_REG_0__SCAN_IN), .A(n3395), .ZN(
        n3394) );
  CLKBUF_X1 U3424 ( .A(n5031), .Z(n5230) );
  NAND2_X1 U3425 ( .A1(n5015), .A2(n5014), .ZN(n5013) );
  NAND2_X1 U3426 ( .A1(n3495), .A2(n3494), .ZN(n4595) );
  CLKBUF_X1 U3427 ( .A(n5191), .Z(n6011) );
  NAND2_X1 U3428 ( .A1(n4602), .A2(n3969), .ZN(n5978) );
  NAND2_X2 U3429 ( .A1(n5421), .A2(n4248), .ZN(n5862) );
  INV_X2 U3430 ( .A(n5537), .ZN(n2945) );
  INV_X2 U3431 ( .A(n6082), .ZN(n6073) );
  AND2_X2 U3432 ( .A1(n4292), .A2(n5190), .ZN(n4247) );
  NAND2_X1 U3433 ( .A1(n4047), .A2(n5190), .ZN(n4691) );
  INV_X1 U3434 ( .A(n4262), .ZN(n4065) );
  INV_X1 U3435 ( .A(n4465), .ZN(n4299) );
  INV_X4 U3436 ( .A(n4275), .ZN(n5190) );
  AND4_X1 U3437 ( .A1(n3134), .A2(n3133), .A3(n3132), .A4(n3131), .ZN(n3140)
         );
  AND4_X1 U3438 ( .A1(n3130), .A2(n3129), .A3(n3128), .A4(n3127), .ZN(n3141)
         );
  AND4_X1 U3439 ( .A1(n2977), .A2(n2976), .A3(n2975), .A4(n2974), .ZN(n2988)
         );
  AND4_X1 U3440 ( .A1(n2973), .A2(n2972), .A3(n2971), .A4(n2970), .ZN(n2989)
         );
  CLKBUF_X3 U3441 ( .A(n2994), .Z(n3941) );
  INV_X2 U3442 ( .A(n5591), .ZN(n2946) );
  AND2_X2 U3443 ( .A1(n5157), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n2959)
         );
  NOR2_X1 U3444 ( .A1(n5157), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n2961)
         );
  AND2_X2 U34450 ( .A1(n5404), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5400) );
  INV_X2 U34460 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6405) );
  NAND4_X1 U34480 ( .A1(n2989), .A2(n2988), .A3(n2987), .A4(n2986), .ZN(n2948)
         );
  NAND4_X1 U3449 ( .A1(n2989), .A2(n2988), .A3(n2987), .A4(n2986), .ZN(n4465)
         );
  AND2_X1 U3450 ( .A1(n3153), .A2(n4116), .ZN(n3261) );
  NAND2_X1 U34510 ( .A1(n4236), .A2(n4275), .ZN(n3153) );
  CLKBUF_X1 U34520 ( .A(n3313), .Z(n3940) );
  CLKBUF_X2 U34530 ( .A(n3312), .Z(n3716) );
  NAND2_X1 U34550 ( .A1(n3490), .A2(n3489), .ZN(n4388) );
  NOR2_X1 U34560 ( .A1(n4247), .A2(n3501), .ZN(n3269) );
  XNOR2_X1 U3457 ( .A(n3326), .B(n3325), .ZN(n3447) );
  AND2_X1 U3458 ( .A1(n2949), .A2(n4960), .ZN(n4944) );
  NOR2_X1 U34590 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n2962) );
  NOR2_X1 U34600 ( .A1(n4719), .A2(n4720), .ZN(n4721) );
  NOR2_X1 U34610 ( .A1(n4116), .A2(n6405), .ZN(n3669) );
  AND2_X1 U34620 ( .A1(n5581), .A2(n5579), .ZN(n5251) );
  OR2_X1 U34630 ( .A1(n4121), .A2(n3100), .ZN(n3055) );
  NAND2_X1 U34640 ( .A1(n3264), .A2(n3263), .ZN(n4011) );
  INV_X1 U34650 ( .A(n4109), .ZN(n4239) );
  OR2_X1 U3466 ( .A1(n3345), .A2(n3344), .ZN(n4696) );
  NAND2_X1 U34680 ( .A1(n5696), .A2(n3448), .ZN(n3427) );
  AND2_X1 U34690 ( .A1(n4072), .A2(n4042), .ZN(n4196) );
  AND4_X1 U34700 ( .A1(n2981), .A2(n2980), .A3(n2979), .A4(n2978), .ZN(n2987)
         );
  OR2_X1 U34710 ( .A1(n5808), .A2(READY_N), .ZN(n4020) );
  INV_X1 U34720 ( .A(n3956), .ZN(n4238) );
  OR2_X1 U34730 ( .A1(n5264), .A2(n5257), .ZN(n5266) );
  NOR2_X2 U34740 ( .A1(n4983), .A2(n4982), .ZN(n5015) );
  INV_X1 U3475 ( .A(n4259), .ZN(n3495) );
  NOR2_X1 U3476 ( .A1(n4260), .A2(n4252), .ZN(n3494) );
  INV_X1 U3477 ( .A(n3441), .ZN(n3453) );
  NAND2_X1 U3478 ( .A1(n5139), .A2(n4973), .ZN(n4974) );
  OR2_X1 U3479 ( .A1(n4807), .A2(n5002), .ZN(n4808) );
  NAND2_X1 U3480 ( .A1(n4196), .A2(n4077), .ZN(n5074) );
  NAND2_X1 U3481 ( .A1(n3305), .A2(n3304), .ZN(n3307) );
  NAND2_X2 U3482 ( .A1(n3235), .A2(n3234), .ZN(n4107) );
  NOR2_X1 U3483 ( .A1(n6255), .A2(n4554), .ZN(n4560) );
  AND4_X1 U3484 ( .A1(n3157), .A2(n3156), .A3(n3155), .A4(n3154), .ZN(n3174)
         );
  AND4_X1 U3485 ( .A1(n3166), .A2(n3165), .A3(n3164), .A4(n3163), .ZN(n3172)
         );
  AND4_X1 U3486 ( .A1(n3161), .A2(n3160), .A3(n3159), .A4(n3158), .ZN(n3173)
         );
  AND4_X1 U3487 ( .A1(n3125), .A2(n3124), .A3(n3123), .A4(n3122), .ZN(n3142)
         );
  NAND2_X1 U3488 ( .A1(n6187), .A2(n4832), .ZN(n6255) );
  INV_X2 U3489 ( .A(n5421), .ZN(n6014) );
  CLKBUF_X1 U3490 ( .A(n4266), .Z(n4554) );
  INV_X1 U3491 ( .A(n5764), .ZN(n5801) );
  NOR2_X1 U3492 ( .A1(n4047), .A2(n3265), .ZN(n3273) );
  AND2_X1 U3493 ( .A1(n4940), .A2(n4939), .ZN(n4941) );
  AND2_X1 U3494 ( .A1(n3260), .A2(n4081), .ZN(n3287) );
  CLKBUF_X2 U3495 ( .A(n3311), .Z(n3930) );
  AOI21_X1 U3496 ( .B1(n6383), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n3194), 
        .ZN(n3195) );
  NOR2_X1 U3497 ( .A1(n3193), .A2(n3197), .ZN(n3194) );
  INV_X1 U3498 ( .A(n3198), .ZN(n3193) );
  AND2_X1 U3499 ( .A1(n3271), .A2(n4280), .ZN(n4001) );
  AND2_X1 U3500 ( .A1(n5453), .A2(n5450), .ZN(n5451) );
  NAND2_X2 U3501 ( .A1(n5477), .A2(n5473), .ZN(n5452) );
  AND2_X1 U3502 ( .A1(n5028), .A2(n5027), .ZN(n5229) );
  OR2_X1 U3503 ( .A1(n5120), .A2(n4945), .ZN(n5037) );
  AND2_X1 U3504 ( .A1(n4959), .A2(n4944), .ZN(n5028) );
  AND2_X1 U3505 ( .A1(n5581), .A2(n6126), .ZN(n4807) );
  OR2_X1 U3506 ( .A1(n3355), .A2(n3354), .ZN(n4354) );
  NAND2_X1 U3507 ( .A1(n3359), .A2(n4692), .ZN(n3385) );
  CLKBUF_X1 U3508 ( .A(n3428), .Z(n3829) );
  OAI21_X1 U3509 ( .B1(n4236), .B2(n4065), .A(n3243), .ZN(n3244) );
  AOI21_X1 U3510 ( .B1(n6520), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n3230), 
        .ZN(n3231) );
  XNOR2_X1 U3511 ( .A(n3447), .B(n3448), .ZN(n4346) );
  INV_X1 U3512 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6372) );
  AND4_X1 U3513 ( .A1(n3170), .A2(n3169), .A3(n3168), .A4(n3167), .ZN(n3171)
         );
  AND4_X1 U3514 ( .A1(n3138), .A2(n3137), .A3(n3136), .A4(n3135), .ZN(n3139)
         );
  AOI21_X1 U3515 ( .B1(n6413), .B2(n4228), .A(n5399), .ZN(n4261) );
  NOR2_X1 U3516 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4261), .ZN(n5708) );
  NAND2_X1 U3517 ( .A1(n3188), .A2(n3187), .ZN(n3987) );
  AND2_X1 U3518 ( .A1(n6503), .A2(n3251), .ZN(n4890) );
  NAND2_X1 U3519 ( .A1(n4154), .A2(n4142), .ZN(n4254) );
  OR2_X1 U3520 ( .A1(n3853), .A2(n3852), .ZN(n3902) );
  AND2_X1 U3521 ( .A1(n5282), .A2(n5178), .ZN(n5210) );
  AND2_X1 U3522 ( .A1(n5282), .A2(n5281), .ZN(n5315) );
  NOR2_X1 U3523 ( .A1(n3890), .A2(n5274), .ZN(n3881) );
  AND2_X1 U3524 ( .A1(n3770), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3891)
         );
  AND2_X1 U3525 ( .A1(n3694), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3695)
         );
  NAND2_X1 U3526 ( .A1(n3695), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3747)
         );
  NOR2_X1 U3527 ( .A1(n3648), .A2(n5166), .ZN(n3675) );
  AND2_X1 U3528 ( .A1(n3675), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3694)
         );
  INV_X1 U3529 ( .A(n5476), .ZN(n5172) );
  NOR2_X1 U3530 ( .A1(n6533), .A2(n3589), .ZN(n3667) );
  INV_X1 U3531 ( .A(n3667), .ZN(n3607) );
  NOR2_X1 U3532 ( .A1(n3574), .A2(n3559), .ZN(n3588) );
  NAND2_X1 U3533 ( .A1(n4721), .A2(n3557), .ZN(n4983) );
  INV_X1 U3534 ( .A(n3525), .ZN(n3526) );
  NAND2_X1 U3535 ( .A1(n4582), .A2(n4581), .ZN(n4719) );
  NOR2_X1 U3536 ( .A1(n3504), .A2(n3503), .ZN(n3505) );
  NAND2_X1 U3537 ( .A1(n3505), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3525)
         );
  AOI21_X1 U3538 ( .B1(n4677), .B2(n3631), .A(n3510), .ZN(n4594) );
  AOI21_X1 U3539 ( .B1(n4388), .B2(n3631), .A(n3493), .ZN(n4252) );
  AOI21_X1 U3540 ( .B1(n4379), .B2(n3631), .A(n3473), .ZN(n4260) );
  NOR2_X1 U3541 ( .A1(n3452), .A2(n4663), .ZN(n3471) );
  AOI21_X1 U3542 ( .B1(n4832), .B2(n3631), .A(n3457), .ZN(n4152) );
  NAND2_X1 U3543 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3441) );
  OR2_X1 U3544 ( .A1(n3405), .A2(n4123), .ZN(n4147) );
  AND2_X1 U3545 ( .A1(n4125), .A2(n4126), .ZN(n4123) );
  NOR2_X1 U3546 ( .A1(n5876), .A2(n5253), .ZN(n5881) );
  NAND2_X1 U3547 ( .A1(n4931), .A2(n3056), .ZN(n5137) );
  OR2_X1 U3548 ( .A1(n4806), .A2(n4925), .ZN(n5002) );
  CLKBUF_X1 U3549 ( .A(n4803), .Z(n5001) );
  AND2_X1 U3550 ( .A1(n3015), .A2(n3014), .ZN(n4070) );
  AND2_X1 U3551 ( .A1(n4074), .A2(n5074), .ZN(n4967) );
  INV_X1 U3552 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4206) );
  INV_X2 U3554 ( .A(n4049), .ZN(n4280) );
  NAND2_X1 U3555 ( .A1(n3413), .A2(n3412), .ZN(n6309) );
  OR2_X1 U3556 ( .A1(n6481), .A2(n4261), .ZN(n4300) );
  AOI21_X1 U3557 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n4761), .A(n5757), .ZN(
        n6259) );
  OR2_X1 U3558 ( .A1(n4890), .A2(n6483), .ZN(n5815) );
  INV_X1 U3559 ( .A(n5815), .ZN(n5991) );
  AND2_X1 U3560 ( .A1(n5418), .A2(n4463), .ZN(n5958) );
  AND2_X1 U3561 ( .A1(n5532), .A2(n4116), .ZN(n5537) );
  INV_X2 U3562 ( .A(n5509), .ZN(n5532) );
  NOR2_X1 U3563 ( .A1(n6014), .A2(n4248), .ZN(n5544) );
  NAND2_X1 U3564 ( .A1(n6058), .A2(n4246), .ZN(n5421) );
  AND2_X1 U3565 ( .A1(n4233), .A2(n4232), .ZN(n4245) );
  AND2_X1 U3566 ( .A1(n4029), .A2(n4028), .ZN(n6020) );
  BUF_X1 U3567 ( .A(n6040), .Z(n6032) );
  INV_X1 U3568 ( .A(n6075), .ZN(n6079) );
  AND2_X1 U3569 ( .A1(n5266), .A2(n5258), .ZN(n5863) );
  INV_X1 U3570 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4663) );
  INV_X1 U3571 ( .A(n6118), .ZN(n5593) );
  AND2_X1 U3572 ( .A1(n5912), .A2(n4131), .ZN(n6109) );
  NAND2_X1 U3573 ( .A1(n4233), .A2(n4127), .ZN(n5912) );
  AND2_X1 U3574 ( .A1(n4077), .A2(n4064), .ZN(n6171) );
  AND2_X1 U3575 ( .A1(n4077), .A2(n6366), .ZN(n4965) );
  INV_X1 U3576 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4761) );
  INV_X1 U3577 ( .A(n6308), .ZN(n6500) );
  INV_X1 U3578 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6376) );
  NAND2_X2 U3579 ( .A1(n4220), .A2(n3310), .ZN(n4894) );
  NAND2_X1 U3580 ( .A1(n3309), .A2(n3308), .ZN(n3310) );
  INV_X1 U3581 ( .A(n4832), .ZN(n6188) );
  CLKBUF_X1 U3582 ( .A(n4523), .Z(n6222) );
  INV_X2 U3583 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5404) );
  INV_X2 U3584 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5157) );
  NOR2_X1 U3585 ( .A1(n4559), .A2(n4766), .ZN(n5764) );
  INV_X1 U3586 ( .A(n5703), .ZN(n5743) );
  NAND2_X1 U3587 ( .A1(n5581), .A2(n4962), .ZN(n2949) );
  NAND2_X1 U3588 ( .A1(n3993), .A2(n3186), .ZN(n4091) );
  INV_X1 U3589 ( .A(n4091), .ZN(n3188) );
  INV_X1 U3590 ( .A(n5282), .ZN(n5264) );
  OR2_X1 U3591 ( .A1(n3985), .A2(n3984), .ZN(U2796) );
  INV_X1 U3592 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5073) );
  OR2_X1 U3593 ( .A1(n3447), .A2(n3427), .ZN(n3496) );
  INV_X1 U3594 ( .A(n3496), .ZN(n3476) );
  NAND2_X1 U3595 ( .A1(n4280), .A2(n3999), .ZN(n4355) );
  INV_X1 U3596 ( .A(n4355), .ZN(n3263) );
  OR2_X1 U3597 ( .A1(n3280), .A2(n3279), .ZN(n2951) );
  NOR2_X1 U3598 ( .A1(n4686), .A2(n6083), .ZN(n2952) );
  AND2_X1 U3599 ( .A1(n3498), .A2(n3497), .ZN(n2953) );
  AND2_X1 U3600 ( .A1(n3219), .A2(n3218), .ZN(n3222) );
  OR2_X1 U3601 ( .A1(n3221), .A2(n3190), .ZN(n3192) );
  INV_X1 U3602 ( .A(n4011), .ZN(n3268) );
  NAND2_X1 U3603 ( .A1(n4236), .A2(n5190), .ZN(n3243) );
  NAND2_X1 U3604 ( .A1(n3192), .A2(n3191), .ZN(n3198) );
  AND2_X1 U3605 ( .A1(n5229), .A2(n5029), .ZN(n5030) );
  NOR2_X1 U3606 ( .A1(n3324), .A2(n3323), .ZN(n4347) );
  NAND2_X1 U3607 ( .A1(n3296), .A2(n3295), .ZN(n3298) );
  AND2_X1 U3608 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4198) );
  AND2_X1 U3609 ( .A1(n4465), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3205) );
  OR2_X1 U3610 ( .A1(n4465), .A2(n6520), .ZN(n3361) );
  INV_X1 U3611 ( .A(n4299), .ZN(n3187) );
  OR2_X1 U3612 ( .A1(n4065), .A2(n6520), .ZN(n4109) );
  AND2_X2 U3613 ( .A1(n4198), .A2(n2962), .ZN(n3935) );
  INV_X1 U3614 ( .A(n3958), .ZN(n3924) );
  INV_X1 U3615 ( .A(n3669), .ZN(n3956) );
  AND2_X1 U3616 ( .A1(n5037), .A2(n5036), .ZN(n5038) );
  NAND2_X1 U3617 ( .A1(n4683), .A2(n4682), .ZN(n4689) );
  AND2_X1 U3618 ( .A1(n4001), .A2(n3272), .ZN(n4235) );
  OR2_X1 U3619 ( .A1(n3991), .A2(n3284), .ZN(n4006) );
  NOR2_X1 U3620 ( .A1(n3501), .A2(n4691), .ZN(n3233) );
  NAND2_X1 U3621 ( .A1(n3381), .A2(n3380), .ZN(n3448) );
  NAND2_X1 U3622 ( .A1(n3205), .A2(n4065), .ZN(n3501) );
  NAND2_X1 U3623 ( .A1(n4109), .A2(n3361), .ZN(n3499) );
  NOR2_X1 U3624 ( .A1(n6183), .A2(n3196), .ZN(n3240) );
  NOR2_X1 U3625 ( .A1(n3902), .A2(n5181), .ZN(n3903) );
  BUF_X1 U3626 ( .A(n3020), .Z(n5078) );
  XNOR2_X1 U3627 ( .A(n4694), .B(n3502), .ZN(n4677) );
  OR2_X1 U3628 ( .A1(n3871), .A2(n5312), .ZN(n3853) );
  AND2_X1 U3629 ( .A1(n5176), .A2(n5175), .ZN(n3751) );
  OR2_X1 U3630 ( .A1(n5013), .A2(n3606), .ZN(n5473) );
  INV_X1 U3631 ( .A(n4920), .ZN(n3557) );
  OR2_X1 U3632 ( .A1(n5252), .A2(n5251), .ZN(n5876) );
  NAND2_X1 U3633 ( .A1(n3476), .A2(n2953), .ZN(n4694) );
  AOI21_X1 U3634 ( .B1(n4406), .B2(n4405), .A(n4365), .ZN(n6111) );
  OR2_X1 U3635 ( .A1(n3328), .A2(n3327), .ZN(n3329) );
  NAND2_X1 U3636 ( .A1(n3232), .A2(n3231), .ZN(n3235) );
  AND2_X1 U3637 ( .A1(n4485), .A2(n4486), .ZN(n4620) );
  OR2_X1 U3638 ( .A1(n3185), .A2(n3184), .ZN(n4049) );
  NAND2_X1 U3639 ( .A1(n4523), .A2(n6520), .ZN(n3426) );
  AOI21_X1 U3640 ( .B1(n3981), .B2(REIP_REG_31__SCAN_IN), .A(n3980), .ZN(n3982) );
  OR2_X1 U3641 ( .A1(n5814), .A2(n3977), .ZN(n5384) );
  NOR2_X1 U3642 ( .A1(n3747), .A2(n5445), .ZN(n3713) );
  NOR2_X1 U3643 ( .A1(n4890), .A2(n6405), .ZN(n4602) );
  NOR2_X1 U3644 ( .A1(n6566), .A2(n3607), .ZN(n3665) );
  NOR2_X1 U3645 ( .A1(n3542), .A2(n3527), .ZN(n3558) );
  OR2_X1 U3646 ( .A1(n3965), .A2(n5379), .ZN(n3967) );
  INV_X1 U3647 ( .A(n4890), .ZN(n4992) );
  AND2_X1 U3648 ( .A1(n4671), .A2(n3048), .ZN(n4931) );
  NAND2_X1 U3649 ( .A1(n3100), .A2(n5078), .ZN(n4068) );
  AND4_X1 U3650 ( .A1(n2985), .A2(n2984), .A3(n2983), .A4(n2982), .ZN(n2986)
         );
  AND2_X1 U3651 ( .A1(n5502), .A2(n5375), .ZN(n5426) );
  AND2_X1 U3652 ( .A1(n3713), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3770)
         );
  AND2_X1 U3653 ( .A1(n5452), .A2(n5474), .ZN(n5476) );
  AND2_X1 U3654 ( .A1(n4262), .A2(n5190), .ZN(n4008) );
  NAND2_X1 U3655 ( .A1(n5047), .A2(n5046), .ZN(n5414) );
  AND2_X1 U3656 ( .A1(n5232), .A2(n5231), .ZN(n5577) );
  AND2_X1 U3657 ( .A1(n5004), .A2(n4810), .ZN(n4940) );
  NAND2_X1 U3658 ( .A1(n4060), .A2(n4059), .ZN(n4077) );
  AND2_X1 U3659 ( .A1(n4100), .A2(n4099), .ZN(n6375) );
  OR2_X1 U3660 ( .A1(n4767), .A2(n4615), .ZN(n4791) );
  INV_X1 U3661 ( .A(n5696), .ZN(n4486) );
  INV_X1 U3662 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6383) );
  NAND2_X1 U3663 ( .A1(n4012), .A2(n4233), .ZN(n5808) );
  OAI21_X1 U3664 ( .B1(n3983), .B2(n5820), .A(n3982), .ZN(n3984) );
  NAND2_X1 U3665 ( .A1(n3891), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3890)
         );
  NAND2_X1 U3666 ( .A1(n3526), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3542)
         );
  INV_X1 U3667 ( .A(n5820), .ZN(n5976) );
  INV_X1 U3668 ( .A(n5983), .ZN(n5992) );
  OAI21_X1 U3669 ( .B1(n5434), .B2(n5359), .A(n5360), .ZN(n3111) );
  NOR2_X1 U3670 ( .A1(n5497), .A2(n3089), .ZN(n5092) );
  NOR2_X1 U3671 ( .A1(n5172), .A2(n5173), .ZN(n5171) );
  INV_X1 U3672 ( .A(n4931), .ZN(n4986) );
  NAND2_X1 U3673 ( .A1(n4256), .A2(n4251), .ZN(n4669) );
  AND2_X1 U3674 ( .A1(n4115), .A2(n4114), .ZN(n5509) );
  NOR2_X1 U3675 ( .A1(n6501), .A2(n6020), .ZN(n6040) );
  OR2_X1 U3676 ( .A1(n4020), .A2(n4284), .ZN(n6058) );
  NOR2_X1 U3677 ( .A1(n5315), .A2(n5285), .ZN(n5829) );
  NOR2_X1 U3678 ( .A1(n5524), .A2(n5523), .ZN(n6008) );
  NAND2_X1 U3679 ( .A1(n5119), .A2(n5118), .ZN(n5477) );
  INV_X1 U3680 ( .A(n4721), .ZN(n4921) );
  NAND2_X1 U3681 ( .A1(n3471), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3504)
         );
  NAND2_X1 U3682 ( .A1(n3453), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3452)
         );
  AND2_X1 U3683 ( .A1(n4107), .A2(n4053), .ZN(n4233) );
  NAND2_X1 U3684 ( .A1(n5414), .A2(n5089), .ZN(n5549) );
  AND2_X1 U3685 ( .A1(n5233), .A2(n5577), .ZN(n5252) );
  OR2_X1 U3686 ( .A1(n4823), .A2(n4965), .ZN(n5052) );
  AND2_X1 U3687 ( .A1(n5052), .A2(n5686), .ZN(n6174) );
  INV_X1 U3688 ( .A(n5708), .ZN(n5757) );
  AND2_X1 U3689 ( .A1(n4107), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5399) );
  INV_X1 U3690 ( .A(n4871), .ZN(n6212) );
  AND2_X1 U3691 ( .A1(n4554), .A2(n4766), .ZN(n6184) );
  INV_X1 U3692 ( .A(n4614), .ZN(n6187) );
  INV_X1 U3693 ( .A(n4791), .ZN(n4649) );
  INV_X1 U3694 ( .A(n4484), .ZN(n4519) );
  INV_X1 U3695 ( .A(n4754), .ZN(n4577) );
  OR2_X1 U3696 ( .A1(n6314), .A2(n6313), .ZN(n6361) );
  AND2_X1 U3697 ( .A1(n4322), .A2(n4615), .ZN(n6359) );
  INV_X1 U3698 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6520) );
  AND2_X1 U3699 ( .A1(n5808), .A2(n5810), .ZN(n6503) );
  OR2_X1 U3700 ( .A1(n5418), .A2(n4462), .ZN(n5820) );
  OR2_X1 U3701 ( .A1(n5210), .A2(n5209), .ZN(n5821) );
  NAND2_X1 U3702 ( .A1(n5264), .A2(n5214), .ZN(n5304) );
  INV_X1 U3703 ( .A(n5544), .ZN(n5127) );
  INV_X1 U3704 ( .A(n6020), .ZN(n6043) );
  NAND2_X1 U3705 ( .A1(n4019), .A2(n4233), .ZN(n6075) );
  OAI21_X1 U3706 ( .B1(n5210), .B2(n5180), .A(n5427), .ZN(n5487) );
  INV_X1 U3707 ( .A(n5829), .ZN(n5310) );
  OR2_X1 U3708 ( .A1(n6109), .A2(n4407), .ZN(n6118) );
  INV_X1 U3709 ( .A(n6171), .ZN(n5680) );
  AND2_X1 U3710 ( .A1(n5712), .A2(n5711), .ZN(n5750) );
  NOR2_X1 U3711 ( .A1(n5759), .A2(n5758), .ZN(n5807) );
  OR2_X1 U3712 ( .A1(n6255), .A2(n4831), .ZN(n6297) );
  OR2_X1 U3713 ( .A1(n6255), .A2(n6252), .ZN(n6364) );
  NOR2_X4 U3714 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5391) );
  NOR2_X4 U3715 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n2963) );
  AOI22_X1 U3716 ( .A1(n3311), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3126), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n2958) );
  AND2_X2 U3717 ( .A1(n2959), .A2(n5400), .ZN(n3337) );
  AND2_X4 U3719 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5152) );
  AND2_X2 U3720 ( .A1(n2961), .A2(n5152), .ZN(n3362) );
  AOI22_X1 U3721 ( .A1(n3337), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n2957) );
  AND2_X2 U3722 ( .A1(n6369), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n2960)
         );
  AND2_X2 U3723 ( .A1(n2960), .A2(n2963), .ZN(n3313) );
  AOI22_X1 U3724 ( .A1(n3312), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n2956) );
  AND2_X2 U3725 ( .A1(n5400), .A2(n4219), .ZN(n3338) );
  AOI22_X1 U3726 ( .A1(n3331), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3338), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n2955) );
  NAND4_X1 U3727 ( .A1(n2958), .A2(n2957), .A3(n2956), .A4(n2955), .ZN(n2969)
         );
  AND2_X2 U3728 ( .A1(n2959), .A2(n5391), .ZN(n3318) );
  AND2_X2 U3729 ( .A1(n2960), .A2(n4219), .ZN(n2994) );
  BUF_X2 U3730 ( .A(n2994), .Z(n3842) );
  AOI22_X1 U3731 ( .A1(n3318), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3842), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n2967) );
  AND2_X2 U3732 ( .A1(n2961), .A2(n5400), .ZN(n3339) );
  AOI22_X1 U3733 ( .A1(n3339), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3935), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n2966) );
  AND2_X2 U3734 ( .A1(n5391), .A2(n2963), .ZN(n3332) );
  AND2_X2 U3735 ( .A1(n2963), .A2(n5152), .ZN(n3162) );
  BUF_X4 U3736 ( .A(n3162), .Z(n3943) );
  AOI22_X1 U3737 ( .A1(n3332), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n2965) );
  AND2_X2 U3738 ( .A1(n5391), .A2(n4219), .ZN(n3179) );
  CLKBUF_X3 U3739 ( .A(n3179), .Z(n3944) );
  AND2_X2 U3740 ( .A1(n4219), .A2(n5152), .ZN(n3428) );
  AOI22_X1 U3741 ( .A1(n3944), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n2964) );
  NAND4_X1 U3742 ( .A1(n2967), .A2(n2966), .A3(n2965), .A4(n2964), .ZN(n2968)
         );
  OR2_X2 U3743 ( .A1(n2969), .A2(n2968), .ZN(n3999) );
  INV_X2 U3744 ( .A(n3999), .ZN(n4288) );
  NAND2_X1 U3745 ( .A1(n3318), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n2973) );
  NAND2_X1 U3746 ( .A1(n3312), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n2972)
         );
  NAND2_X1 U3747 ( .A1(n3311), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n2971) );
  NAND2_X1 U3748 ( .A1(n3338), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n2970)
         );
  NAND2_X1 U3749 ( .A1(n3331), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n2977)
         );
  NAND2_X1 U3750 ( .A1(n3337), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n2976) );
  NAND2_X1 U3751 ( .A1(n3313), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n2975) );
  NAND2_X1 U3752 ( .A1(n3126), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n2974) );
  NAND2_X1 U3753 ( .A1(n3362), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n2981) );
  NAND2_X1 U3754 ( .A1(n3941), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n2980)
         );
  NAND2_X1 U3755 ( .A1(n3428), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n2979)
         );
  NAND2_X1 U3756 ( .A1(n3823), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n2978) );
  NAND2_X1 U3757 ( .A1(n3339), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n2985) );
  NAND2_X1 U3758 ( .A1(n3332), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n2984) );
  NAND2_X1 U3759 ( .A1(n3732), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n2983)
         );
  NAND2_X1 U3760 ( .A1(n3935), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n2982) );
  AOI22_X1 U3761 ( .A1(n3312), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n2993) );
  AOI22_X1 U3762 ( .A1(n3337), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3338), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n2992) );
  AOI22_X1 U3763 ( .A1(n3331), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n2991) );
  AOI22_X1 U3764 ( .A1(n3126), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n2990) );
  NAND4_X1 U3765 ( .A1(n2993), .A2(n2992), .A3(n2991), .A4(n2990), .ZN(n3000)
         );
  BUF_X2 U3766 ( .A(n2994), .Z(n3915) );
  AOI22_X1 U3767 ( .A1(n3915), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n2998) );
  AOI22_X1 U3768 ( .A1(n3318), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3732), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n2997) );
  AOI22_X1 U3769 ( .A1(n3311), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n2996) );
  AOI22_X1 U3770 ( .A1(n3339), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3935), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n2995) );
  NAND4_X1 U3771 ( .A1(n2998), .A2(n2997), .A3(n2996), .A4(n2995), .ZN(n2999)
         );
  OR2_X4 U3772 ( .A1(n3000), .A2(n2999), .ZN(n4047) );
  NAND2_X1 U3773 ( .A1(n3999), .A2(n4047), .ZN(n3020) );
  NAND2_X1 U3774 ( .A1(n4068), .A2(EBX_REG_16__SCAN_IN), .ZN(n3002) );
  NAND2_X1 U3775 ( .A1(n4047), .A2(n2948), .ZN(n3004) );
  NAND2_X1 U3776 ( .A1(n4092), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3001) );
  NAND2_X1 U3777 ( .A1(n3002), .A2(n3001), .ZN(n3003) );
  XNOR2_X1 U3778 ( .A(n3003), .B(n5078), .ZN(n5146) );
  INV_X2 U3779 ( .A(n3004), .ZN(n4121) );
  NAND2_X1 U3780 ( .A1(n4121), .A2(n5078), .ZN(n3097) );
  NAND2_X1 U3781 ( .A1(n5078), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3005) );
  OAI211_X1 U3782 ( .C1(n4092), .C2(EBX_REG_13__SCAN_IN), .A(n3100), .B(n3005), 
        .ZN(n3006) );
  OAI21_X1 U3783 ( .B1(n3097), .B2(EBX_REG_13__SCAN_IN), .A(n3006), .ZN(n5138)
         );
  INV_X2 U3784 ( .A(n3020), .ZN(n5432) );
  NAND2_X1 U3785 ( .A1(n5432), .A2(EBX_REG_5__SCAN_IN), .ZN(n3009) );
  INV_X1 U3786 ( .A(n3097), .ZN(n3082) );
  INV_X1 U3787 ( .A(EBX_REG_5__SCAN_IN), .ZN(n3007) );
  NAND2_X1 U3788 ( .A1(n3082), .A2(n3007), .ZN(n3008) );
  OAI211_X1 U3789 ( .C1(n4068), .C2(INSTADDRPOINTER_REG_5__SCAN_IN), .A(n3009), 
        .B(n3008), .ZN(n4255) );
  AND2_X4 U3790 ( .A1(n5432), .A2(n4121), .ZN(n3106) );
  INV_X1 U3791 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3010) );
  NAND2_X1 U3792 ( .A1(n3106), .A2(n3010), .ZN(n3013) );
  OR2_X1 U3793 ( .A1(n3100), .A2(n3010), .ZN(n3012) );
  INV_X1 U3794 ( .A(n4121), .ZN(n3064) );
  NAND3_X1 U3795 ( .A1(n3020), .A2(n3064), .A3(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n3011) );
  NAND4_X1 U3796 ( .A1(n3055), .A2(n3013), .A3(n3012), .A4(n3011), .ZN(n3016)
         );
  INV_X1 U3797 ( .A(n3016), .ZN(n3018) );
  NAND2_X1 U3798 ( .A1(n3100), .A2(EBX_REG_0__SCAN_IN), .ZN(n3015) );
  INV_X1 U3799 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4120) );
  NAND2_X1 U3800 ( .A1(n3020), .A2(n4120), .ZN(n3014) );
  XNOR2_X1 U3801 ( .A(n3016), .B(n4070), .ZN(n4122) );
  NOR2_X1 U3802 ( .A1(n4122), .A2(n4092), .ZN(n3017) );
  NOR2_X1 U3803 ( .A1(n3018), .A2(n3017), .ZN(n4149) );
  INV_X1 U3804 ( .A(EBX_REG_2__SCAN_IN), .ZN(n3019) );
  NAND2_X1 U3805 ( .A1(n3106), .A2(n3019), .ZN(n3024) );
  INV_X1 U3806 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U3807 ( .A1(n3100), .A2(n6173), .ZN(n3022) );
  NAND2_X1 U3808 ( .A1(n4121), .A2(n3019), .ZN(n3021) );
  NAND3_X1 U3809 ( .A1(n3022), .A2(n3021), .A3(n5078), .ZN(n3023) );
  NAND2_X1 U3810 ( .A1(n3024), .A2(n3023), .ZN(n4150) );
  NAND2_X1 U3811 ( .A1(n4149), .A2(n4150), .ZN(n4155) );
  NAND2_X1 U3812 ( .A1(n5078), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3025)
         );
  OAI211_X1 U3813 ( .C1(n4092), .C2(EBX_REG_3__SCAN_IN), .A(n3100), .B(n3025), 
        .ZN(n3026) );
  OAI21_X1 U3814 ( .B1(n3097), .B2(EBX_REG_3__SCAN_IN), .A(n3026), .ZN(n4156)
         );
  NOR2_X2 U3815 ( .A1(n4155), .A2(n4156), .ZN(n4154) );
  INV_X1 U3816 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6594) );
  NAND2_X1 U3817 ( .A1(n3106), .A2(n6594), .ZN(n3030) );
  INV_X1 U3818 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6159) );
  NAND2_X1 U3819 ( .A1(n3100), .A2(n6159), .ZN(n3028) );
  NAND2_X1 U3820 ( .A1(n4121), .A2(n6594), .ZN(n3027) );
  NAND3_X1 U3821 ( .A1(n3028), .A2(n3027), .A3(n5078), .ZN(n3029) );
  NAND2_X1 U3822 ( .A1(n3030), .A2(n3029), .ZN(n4142) );
  NOR2_X2 U3823 ( .A1(n4255), .A2(n4254), .ZN(n4256) );
  INV_X1 U3824 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4469) );
  NAND2_X1 U3825 ( .A1(n3106), .A2(n4469), .ZN(n3033) );
  OR2_X1 U3826 ( .A1(n3100), .A2(n4469), .ZN(n3032) );
  NAND2_X1 U3827 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4092), .ZN(n3031)
         );
  NAND4_X1 U3828 ( .A1(n3055), .A2(n3033), .A3(n3032), .A4(n3031), .ZN(n4251)
         );
  NAND2_X1 U3829 ( .A1(n5432), .A2(EBX_REG_7__SCAN_IN), .ZN(n3035) );
  OR2_X1 U3830 ( .A1(n4068), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3034)
         );
  OAI211_X1 U3831 ( .C1(EBX_REG_7__SCAN_IN), .C2(n3097), .A(n3035), .B(n3034), 
        .ZN(n4670) );
  NOR2_X2 U3832 ( .A1(n4669), .A2(n4670), .ZN(n4671) );
  INV_X1 U3833 ( .A(EBX_REG_10__SCAN_IN), .ZN(n3036) );
  NAND2_X1 U3834 ( .A1(n3106), .A2(n3036), .ZN(n3039) );
  OR2_X1 U3835 ( .A1(n3100), .A2(n3036), .ZN(n3038) );
  NAND2_X1 U3836 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n4092), .ZN(n3037) );
  NAND4_X1 U3837 ( .A1(n3055), .A2(n3039), .A3(n3038), .A4(n3037), .ZN(n4933)
         );
  INV_X1 U3838 ( .A(n4933), .ZN(n3042) );
  NAND2_X1 U3839 ( .A1(n5432), .A2(EBX_REG_9__SCAN_IN), .ZN(n3041) );
  INV_X1 U3840 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4880) );
  NAND2_X1 U3841 ( .A1(n3082), .A2(n4880), .ZN(n3040) );
  OAI211_X1 U3842 ( .C1(n4068), .C2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n3041), 
        .B(n3040), .ZN(n4879) );
  NOR2_X1 U3843 ( .A1(n3042), .A2(n4879), .ZN(n3047) );
  INV_X1 U3844 ( .A(EBX_REG_8__SCAN_IN), .ZN(n3043) );
  NAND2_X1 U3845 ( .A1(n3106), .A2(n3043), .ZN(n3046) );
  OR2_X1 U3846 ( .A1(n3100), .A2(n3043), .ZN(n3045) );
  NAND2_X1 U3847 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n4092), .ZN(n3044)
         );
  NAND4_X1 U3848 ( .A1(n3055), .A2(n3046), .A3(n3045), .A4(n3044), .ZN(n4584)
         );
  AND2_X1 U3849 ( .A1(n3047), .A2(n4584), .ZN(n3048) );
  INV_X1 U3850 ( .A(EBX_REG_11__SCAN_IN), .ZN(n3051) );
  INV_X1 U3851 ( .A(n4068), .ZN(n3049) );
  INV_X1 U3852 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6126) );
  AOI22_X1 U3853 ( .A1(n3049), .A2(n6126), .B1(n3082), .B2(n3051), .ZN(n3050)
         );
  OAI21_X1 U3854 ( .B1(n5078), .B2(n3051), .A(n3050), .ZN(n4987) );
  INV_X1 U3855 ( .A(n4987), .ZN(n4821) );
  INV_X1 U3856 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5020) );
  NAND2_X1 U3857 ( .A1(n3106), .A2(n5020), .ZN(n3054) );
  OR2_X1 U3858 ( .A1(n3100), .A2(n5020), .ZN(n3053) );
  NAND2_X1 U3859 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n4092), .ZN(n3052) );
  NAND4_X1 U3860 ( .A1(n3055), .A2(n3054), .A3(n3053), .A4(n3052), .ZN(n4822)
         );
  AND2_X1 U3861 ( .A1(n4821), .A2(n4822), .ZN(n3056) );
  NOR2_X2 U3862 ( .A1(n5138), .A2(n5137), .ZN(n5139) );
  INV_X1 U3863 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U3864 ( .A1(n3106), .A2(n5533), .ZN(n3060) );
  INV_X1 U3865 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4962) );
  NAND2_X1 U3866 ( .A1(n3100), .A2(n4962), .ZN(n3058) );
  NAND2_X1 U3867 ( .A1(n4121), .A2(n5533), .ZN(n3057) );
  NAND3_X1 U3868 ( .A1(n3058), .A2(n3057), .A3(n5078), .ZN(n3059) );
  NAND2_X1 U3869 ( .A1(n3060), .A2(n3059), .ZN(n4973) );
  NAND2_X1 U3870 ( .A1(n5432), .A2(EBX_REG_15__SCAN_IN), .ZN(n3062) );
  OR2_X1 U3871 ( .A1(n4068), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3061)
         );
  OAI211_X1 U3872 ( .C1(EBX_REG_15__SCAN_IN), .C2(n3097), .A(n3062), .B(n3061), 
        .ZN(n4948) );
  NOR2_X2 U3873 ( .A1(n4974), .A2(n4948), .ZN(n5145) );
  NAND2_X1 U3874 ( .A1(n5146), .A2(n5145), .ZN(n5526) );
  NAND2_X1 U3875 ( .A1(n5078), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3063) );
  OAI211_X1 U3876 ( .C1(n3064), .C2(EBX_REG_17__SCAN_IN), .A(n3100), .B(n3063), 
        .ZN(n3065) );
  OAI21_X1 U3877 ( .B1(n3097), .B2(EBX_REG_17__SCAN_IN), .A(n3065), .ZN(n5525)
         );
  OR2_X2 U3878 ( .A1(n5526), .A2(n5525), .ZN(n5528) );
  INV_X1 U3879 ( .A(n3100), .ZN(n3086) );
  AOI22_X1 U3880 ( .A1(n3086), .A2(EBX_REG_19__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n4092), .ZN(n3067) );
  INV_X1 U3881 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U3882 ( .A1(n3106), .A2(n5517), .ZN(n3066) );
  AND2_X1 U3883 ( .A1(n3067), .A2(n3066), .ZN(n5082) );
  OR2_X2 U3884 ( .A1(n5528), .A2(n5082), .ZN(n5106) );
  OR2_X1 U3885 ( .A1(n4068), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3069)
         );
  INV_X1 U3886 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U3887 ( .A1(n4121), .A2(n5443), .ZN(n3068) );
  AND2_X1 U3888 ( .A1(n3069), .A2(n3068), .ZN(n5107) );
  OR2_X1 U3889 ( .A1(n4068), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3070)
         );
  INV_X1 U3890 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U3891 ( .A1(n4121), .A2(n5457), .ZN(n5079) );
  NAND2_X1 U3892 ( .A1(n3070), .A2(n5079), .ZN(n5105) );
  NAND2_X1 U3893 ( .A1(n5105), .A2(n5078), .ZN(n3072) );
  NAND2_X1 U3894 ( .A1(n5432), .A2(EBX_REG_20__SCAN_IN), .ZN(n3071) );
  OAI211_X1 U3895 ( .C1(n5107), .C2(n5105), .A(n3072), .B(n3071), .ZN(n3073)
         );
  NOR2_X4 U3896 ( .A1(n5106), .A2(n3073), .ZN(n5506) );
  INV_X1 U3897 ( .A(n3106), .ZN(n3094) );
  NAND2_X1 U3898 ( .A1(n4092), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3075) );
  NAND2_X1 U3899 ( .A1(n3086), .A2(EBX_REG_23__SCAN_IN), .ZN(n3074) );
  OAI211_X1 U3900 ( .C1(n3094), .C2(EBX_REG_23__SCAN_IN), .A(n3075), .B(n3074), 
        .ZN(n5494) );
  AOI22_X1 U3901 ( .A1(n3086), .A2(EBX_REG_21__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n4092), .ZN(n3078) );
  INV_X1 U3902 ( .A(EBX_REG_21__SCAN_IN), .ZN(n3076) );
  NAND2_X1 U3903 ( .A1(n3106), .A2(n3076), .ZN(n3077) );
  AND2_X1 U3904 ( .A1(n3078), .A2(n3077), .ZN(n5505) );
  OR2_X1 U3905 ( .A1(n4068), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3080)
         );
  NAND2_X1 U3906 ( .A1(n5432), .A2(EBX_REG_22__SCAN_IN), .ZN(n3079) );
  OAI211_X1 U3907 ( .C1(EBX_REG_22__SCAN_IN), .C2(n3097), .A(n3080), .B(n3079), 
        .ZN(n5218) );
  NOR2_X1 U3908 ( .A1(n5505), .A2(n5218), .ZN(n5217) );
  AND2_X1 U3909 ( .A1(n5494), .A2(n5217), .ZN(n3081) );
  NAND2_X2 U3910 ( .A1(n5506), .A2(n3081), .ZN(n5497) );
  OR2_X1 U3911 ( .A1(n4068), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3085)
         );
  INV_X1 U3912 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U3913 ( .A1(n3082), .A2(n5309), .ZN(n3084) );
  NAND2_X1 U3914 ( .A1(n5432), .A2(EBX_REG_25__SCAN_IN), .ZN(n3083) );
  AND3_X1 U3915 ( .A1(n3085), .A2(n3084), .A3(n3083), .ZN(n5067) );
  NAND2_X1 U3916 ( .A1(n4092), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3088) );
  NAND2_X1 U3917 ( .A1(n3086), .A2(EBX_REG_24__SCAN_IN), .ZN(n3087) );
  OAI211_X1 U3918 ( .C1(n3094), .C2(EBX_REG_24__SCAN_IN), .A(n3088), .B(n3087), 
        .ZN(n5270) );
  NAND2_X1 U3919 ( .A1(n5067), .A2(n5270), .ZN(n3089) );
  INV_X1 U3920 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6581) );
  NAND2_X1 U3921 ( .A1(n3100), .A2(n6581), .ZN(n3092) );
  INV_X1 U3922 ( .A(EBX_REG_26__SCAN_IN), .ZN(n3090) );
  NAND2_X1 U3923 ( .A1(n4121), .A2(n3090), .ZN(n3091) );
  NAND3_X1 U3924 ( .A1(n3092), .A2(n5078), .A3(n3091), .ZN(n3093) );
  OAI21_X1 U3925 ( .B1(n3094), .B2(EBX_REG_26__SCAN_IN), .A(n3093), .ZN(n5091)
         );
  NAND2_X1 U3926 ( .A1(n5092), .A2(n5091), .ZN(n5490) );
  OR2_X1 U3927 ( .A1(n4068), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3096)
         );
  NAND2_X1 U3928 ( .A1(n5432), .A2(EBX_REG_27__SCAN_IN), .ZN(n3095) );
  OAI211_X1 U3929 ( .C1(EBX_REG_27__SCAN_IN), .C2(n3097), .A(n3096), .B(n3095), 
        .ZN(n5489) );
  OR2_X2 U3930 ( .A1(n5490), .A2(n5489), .ZN(n5492) );
  OR2_X1 U3931 ( .A1(n4068), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3099)
         );
  INV_X1 U3932 ( .A(EBX_REG_29__SCAN_IN), .ZN(n3105) );
  NAND2_X1 U3933 ( .A1(n4121), .A2(n3105), .ZN(n3098) );
  NAND2_X1 U3934 ( .A1(n3099), .A2(n3098), .ZN(n5431) );
  INV_X1 U3935 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U3936 ( .A1(n3106), .A2(n5488), .ZN(n3103) );
  INV_X1 U3937 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U3938 ( .A1(n3100), .A2(n5186), .ZN(n3101) );
  OAI211_X1 U3939 ( .C1(EBX_REG_28__SCAN_IN), .C2(n4092), .A(n3101), .B(n5078), 
        .ZN(n3102) );
  AND2_X1 U3940 ( .A1(n3103), .A2(n3102), .ZN(n5195) );
  OR2_X1 U3941 ( .A1(n5431), .A2(n5195), .ZN(n3104) );
  OR2_X2 U3942 ( .A1(n5492), .A2(n5195), .ZN(n5430) );
  NAND2_X1 U3943 ( .A1(n3106), .A2(n3105), .ZN(n5429) );
  NOR2_X1 U3944 ( .A1(n5430), .A2(n5429), .ZN(n3107) );
  AOI21_X1 U3945 ( .B1(n5361), .B2(n5078), .A(n3107), .ZN(n5434) );
  NAND2_X1 U3946 ( .A1(n4068), .A2(EBX_REG_30__SCAN_IN), .ZN(n3109) );
  NAND2_X1 U3947 ( .A1(n4092), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3108) );
  NAND2_X1 U3948 ( .A1(n3109), .A2(n3108), .ZN(n5359) );
  INV_X1 U3949 ( .A(n5361), .ZN(n5357) );
  NAND2_X1 U3950 ( .A1(n5357), .A2(n5078), .ZN(n5360) );
  OAI22_X1 U3951 ( .A1(n4068), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4092), .ZN(n3110) );
  XNOR2_X1 U3952 ( .A(n3111), .B(n3110), .ZN(n5608) );
  AOI22_X1 U3953 ( .A1(n3312), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3337), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3115) );
  AOI22_X1 U3954 ( .A1(n3311), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3114) );
  AOI22_X1 U3955 ( .A1(n3339), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3935), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3113) );
  AOI22_X1 U3956 ( .A1(n3331), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3112) );
  NAND4_X1 U3957 ( .A1(n3115), .A2(n3114), .A3(n3113), .A4(n3112), .ZN(n3121)
         );
  AOI22_X1 U3958 ( .A1(n3318), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3842), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3119) );
  AOI22_X1 U3959 ( .A1(n3338), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3126), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3118) );
  AOI22_X1 U3960 ( .A1(n3313), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3117) );
  AOI22_X1 U3961 ( .A1(n3332), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3162), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3116) );
  NAND4_X1 U3962 ( .A1(n3119), .A2(n3118), .A3(n3117), .A4(n3116), .ZN(n3120)
         );
  OR2_X2 U3963 ( .A1(n3121), .A2(n3120), .ZN(n4236) );
  NAND2_X1 U3964 ( .A1(n3362), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3125) );
  NAND2_X1 U3965 ( .A1(n3337), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3124) );
  NAND2_X1 U3966 ( .A1(n3312), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3123)
         );
  NAND2_X1 U3967 ( .A1(n3313), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3122) );
  NAND2_X1 U3968 ( .A1(n3126), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3130) );
  NAND2_X1 U3969 ( .A1(n3331), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3129)
         );
  NAND2_X1 U3970 ( .A1(n3311), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3128) );
  NAND2_X1 U3971 ( .A1(n3338), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3127)
         );
  NAND2_X1 U3972 ( .A1(n3318), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3134) );
  NAND2_X1 U3973 ( .A1(n3941), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3133)
         );
  NAND2_X1 U3974 ( .A1(n3823), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3132) );
  NAND2_X1 U3975 ( .A1(n3332), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3131) );
  NAND2_X1 U3976 ( .A1(n3339), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3138) );
  NAND2_X1 U3977 ( .A1(n3935), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3137) );
  NAND2_X1 U3978 ( .A1(n3732), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3136)
         );
  NAND2_X1 U3979 ( .A1(n3428), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3135)
         );
  AND4_X2 U3980 ( .A1(n3142), .A2(n3141), .A3(n3140), .A4(n3139), .ZN(n4275)
         );
  AOI22_X1 U3981 ( .A1(n3339), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3146) );
  AOI22_X1 U3982 ( .A1(n3311), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3126), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3145) );
  AOI22_X1 U3983 ( .A1(n3312), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3338), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3144) );
  AOI22_X1 U3984 ( .A1(n3362), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3143) );
  NAND4_X1 U3985 ( .A1(n3146), .A2(n3145), .A3(n3144), .A4(n3143), .ZN(n3152)
         );
  AOI22_X1 U3986 ( .A1(n3331), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3150) );
  AOI22_X1 U3987 ( .A1(n3823), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3935), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3149) );
  AOI22_X1 U3988 ( .A1(n3318), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3148) );
  AOI22_X1 U3989 ( .A1(n3337), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3147) );
  NAND4_X1 U3990 ( .A1(n3150), .A2(n3149), .A3(n3148), .A4(n3147), .ZN(n3151)
         );
  OR2_X2 U3991 ( .A1(n3152), .A2(n3151), .ZN(n4116) );
  NAND2_X1 U3992 ( .A1(n3362), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3157) );
  NAND2_X1 U3993 ( .A1(n3337), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3156) );
  NAND2_X1 U3994 ( .A1(n3312), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3155)
         );
  NAND2_X1 U3995 ( .A1(n3313), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3154) );
  NAND2_X1 U3996 ( .A1(n3126), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3161) );
  NAND2_X1 U3997 ( .A1(n3331), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3160)
         );
  NAND2_X1 U3998 ( .A1(n3311), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3159) );
  NAND2_X1 U3999 ( .A1(n3338), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3158)
         );
  NAND2_X1 U4000 ( .A1(n3318), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3166) );
  NAND2_X1 U4001 ( .A1(n3941), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3165)
         );
  NAND2_X1 U4002 ( .A1(n3162), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3164) );
  NAND2_X1 U4003 ( .A1(n3332), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3163) );
  NAND2_X1 U4004 ( .A1(n3339), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3170) );
  NAND2_X1 U4005 ( .A1(n3935), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3169) );
  NAND2_X1 U4006 ( .A1(n3732), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3168)
         );
  NAND2_X1 U4007 ( .A1(n3428), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3167)
         );
  NAND2_X1 U4009 ( .A1(n3261), .A2(n4262), .ZN(n3259) );
  INV_X2 U4010 ( .A(n4236), .ZN(n4292) );
  NOR2_X2 U4011 ( .A1(n3259), .A2(n4247), .ZN(n3993) );
  AOI22_X1 U4012 ( .A1(n3337), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3178) );
  AOI22_X1 U4013 ( .A1(n3312), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3177) );
  AOI22_X1 U4014 ( .A1(n3318), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3338), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3176) );
  AOI22_X1 U4015 ( .A1(n3332), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3175) );
  NAND4_X1 U4016 ( .A1(n3178), .A2(n3177), .A3(n3176), .A4(n3175), .ZN(n3185)
         );
  AOI22_X1 U4017 ( .A1(n3362), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3126), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3183) );
  AOI22_X1 U4018 ( .A1(n3941), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3182) );
  AOI22_X1 U4019 ( .A1(n3339), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3935), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U4020 ( .A1(n3331), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3180) );
  NAND4_X1 U4021 ( .A1(n3183), .A2(n3182), .A3(n3181), .A4(n3180), .ZN(n3184)
         );
  NOR2_X1 U4022 ( .A1(n4355), .A2(n4236), .ZN(n3186) );
  INV_X1 U4023 ( .A(n3987), .ZN(n4012) );
  INV_X1 U4024 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6607) );
  NAND2_X1 U4025 ( .A1(n4761), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3204) );
  INV_X1 U4026 ( .A(n3204), .ZN(n3189) );
  XNOR2_X1 U4027 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3201) );
  AOI22_X1 U4028 ( .A1(n3189), .A2(n3201), .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n6372), .ZN(n3221) );
  XNOR2_X1 U4029 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3220) );
  INV_X1 U4030 ( .A(n3220), .ZN(n3190) );
  NAND2_X1 U4031 ( .A1(n6376), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3191) );
  XNOR2_X1 U4032 ( .A(n4206), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3197)
         );
  OAI222_X1 U4033 ( .A1(n6607), .A2(n3195), .B1(n6607), .B2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C1(n3195), .C2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3236) );
  NAND2_X1 U4034 ( .A1(n3236), .A2(n3499), .ZN(n3232) );
  INV_X1 U4035 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U4036 ( .A1(n3195), .A2(n6607), .ZN(n3196) );
  XNOR2_X1 U4037 ( .A(n3198), .B(n3197), .ZN(n3239) );
  INV_X1 U4038 ( .A(n3239), .ZN(n3199) );
  OAI21_X1 U4039 ( .B1(n3240), .B2(n3199), .A(n3501), .ZN(n3228) );
  NAND2_X1 U4040 ( .A1(n4275), .A2(n3187), .ZN(n3200) );
  NAND2_X1 U4041 ( .A1(n3200), .A2(n4284), .ZN(n3206) );
  INV_X1 U4042 ( .A(n3206), .ZN(n3224) );
  XNOR2_X1 U4043 ( .A(n3201), .B(n3204), .ZN(n3238) );
  NAND2_X1 U4044 ( .A1(n3499), .A2(n4047), .ZN(n3202) );
  NAND2_X1 U4045 ( .A1(n3202), .A2(n5190), .ZN(n3215) );
  NAND2_X1 U4046 ( .A1(n6369), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3203) );
  NAND2_X1 U4047 ( .A1(n3204), .A2(n3203), .ZN(n3208) );
  OAI21_X1 U4048 ( .B1(n4008), .B2(n3208), .A(n3205), .ZN(n3207) );
  NAND2_X1 U4049 ( .A1(n3207), .A2(n3206), .ZN(n3214) );
  INV_X1 U4050 ( .A(n3499), .ZN(n3209) );
  NOR2_X1 U4051 ( .A1(n3209), .A2(n3208), .ZN(n3210) );
  OAI211_X1 U4052 ( .C1(n3238), .C2(n3215), .A(n3214), .B(n3210), .ZN(n3213)
         );
  INV_X1 U4053 ( .A(n3233), .ZN(n3212) );
  NAND3_X1 U4054 ( .A1(n3215), .A2(STATE2_REG_0__SCAN_IN), .A3(n3238), .ZN(
        n3211) );
  NAND3_X1 U4055 ( .A1(n3213), .A2(n3212), .A3(n3211), .ZN(n3219) );
  INV_X1 U4056 ( .A(n3214), .ZN(n3217) );
  INV_X1 U4057 ( .A(n3215), .ZN(n3216) );
  NAND3_X1 U4058 ( .A1(n3217), .A2(n3216), .A3(n3238), .ZN(n3218) );
  XNOR2_X1 U4059 ( .A(n3221), .B(n3220), .ZN(n3237) );
  OAI211_X1 U4060 ( .C1(n3224), .C2(n3222), .A(n3237), .B(n3499), .ZN(n3226)
         );
  NOR2_X1 U4061 ( .A1(n3237), .A2(n3501), .ZN(n3223) );
  OAI21_X1 U4062 ( .B1(n3224), .B2(n3223), .A(n3222), .ZN(n3225) );
  OAI211_X1 U4063 ( .C1(n3239), .C2(n4691), .A(n3226), .B(n3225), .ZN(n3227)
         );
  AOI22_X1 U4064 ( .A1(n3233), .A2(n3240), .B1(n3228), .B2(n3227), .ZN(n3229)
         );
  INV_X1 U4065 ( .A(n3229), .ZN(n3230) );
  NAND2_X1 U4066 ( .A1(n3236), .A2(n3233), .ZN(n3234) );
  INV_X1 U4067 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4237) );
  AND2_X1 U4068 ( .A1(n4237), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3410) );
  NAND2_X1 U4069 ( .A1(n3410), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6407) );
  INV_X1 U4070 ( .A(n6407), .ZN(n4053) );
  INV_X1 U4071 ( .A(n3236), .ZN(n3242) );
  NAND3_X1 U4072 ( .A1(n3239), .A2(n3238), .A3(n3237), .ZN(n3241) );
  AOI21_X1 U4073 ( .B1(n3242), .B2(n3241), .A(n3240), .ZN(n4048) );
  NAND2_X1 U4074 ( .A1(n3244), .A2(n4280), .ZN(n3245) );
  OAI211_X1 U4075 ( .C1(n4247), .C2(n4288), .A(n3245), .B(n4116), .ZN(n3258)
         );
  NAND3_X1 U4076 ( .A1(n4008), .A2(n4299), .A3(n4236), .ZN(n3246) );
  NOR2_X2 U4077 ( .A1(n3258), .A2(n3246), .ZN(n4026) );
  NAND2_X1 U4078 ( .A1(n4026), .A2(n4053), .ZN(n3247) );
  OR2_X1 U4079 ( .A1(n4048), .A2(n3247), .ZN(n5810) );
  INV_X1 U4080 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U4081 ( .A1(n4237), .A2(n6405), .ZN(n6413) );
  NOR3_X1 U4082 ( .A1(n6483), .A2(n6520), .A3(n6413), .ZN(n6400) );
  AND2_X1 U4083 ( .A1(n6520), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3248) );
  NOR2_X1 U4084 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3650) );
  AND2_X1 U4085 ( .A1(n3248), .A2(n3650), .ZN(n6409) );
  INV_X1 U4086 ( .A(n6409), .ZN(n3249) );
  NOR2_X1 U4087 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n5900) );
  NAND2_X1 U4088 ( .A1(n5900), .A2(n6520), .ZN(n4129) );
  OR2_X1 U4089 ( .A1(n4129), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U4090 ( .A1(n3249), .A2(n5585), .ZN(n3250) );
  NOR2_X1 U4091 ( .A1(n6400), .A2(n3250), .ZN(n3251) );
  NOR2_X1 U4092 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3968) );
  INV_X1 U4093 ( .A(n3968), .ZN(n4464) );
  NAND2_X1 U4094 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4464), .ZN(n3252) );
  NOR2_X1 U4095 ( .A1(n4092), .A2(n3252), .ZN(n3253) );
  NAND2_X1 U4096 ( .A1(n4602), .A2(n3253), .ZN(n5983) );
  NAND2_X1 U4097 ( .A1(n5991), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3255)
         );
  AND2_X2 U4098 ( .A1(n4284), .A2(n4465), .ZN(n4697) );
  INV_X1 U4099 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6548) );
  XNOR2_X1 U4100 ( .A(n6548), .B(STATE_REG_1__SCAN_IN), .ZN(n3265) );
  INV_X1 U4101 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6424) );
  NAND2_X1 U4102 ( .A1(n3265), .A2(n6424), .ZN(n6422) );
  INV_X1 U4103 ( .A(n6422), .ZN(n4028) );
  NAND2_X1 U4104 ( .A1(n4028), .A2(n3968), .ZN(n6399) );
  NAND4_X1 U4105 ( .A1(n4602), .A2(n4697), .A3(EBX_REG_31__SCAN_IN), .A4(n6399), .ZN(n3254) );
  OAI211_X1 U4106 ( .C1(n5608), .C2(n5983), .A(n3255), .B(n3254), .ZN(n3985)
         );
  NAND2_X1 U4107 ( .A1(n6405), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3885) );
  INV_X1 U4108 ( .A(n3885), .ZN(n3668) );
  AOI22_X1 U4109 ( .A1(n4238), .A2(EAX_REG_31__SCAN_IN), .B1(n3668), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3964) );
  AOI21_X1 U4110 ( .B1(n4292), .B2(n4049), .A(n4047), .ZN(n3256) );
  OAI21_X1 U4111 ( .B1(n4008), .B2(n4280), .A(n3256), .ZN(n3257) );
  OAI21_X1 U4112 ( .B1(n3258), .B2(n3257), .A(n4299), .ZN(n3286) );
  NAND2_X1 U4113 ( .A1(n3259), .A2(n4697), .ZN(n3260) );
  NAND2_X1 U4114 ( .A1(n4000), .A2(n3999), .ZN(n4081) );
  NAND2_X1 U4115 ( .A1(n4247), .A2(n4262), .ZN(n3262) );
  NAND2_X1 U4116 ( .A1(n3262), .A2(n3261), .ZN(n3995) );
  INV_X1 U4117 ( .A(n3995), .ZN(n3264) );
  INV_X1 U4118 ( .A(n3273), .ZN(n3266) );
  NAND2_X1 U4119 ( .A1(n3266), .A2(n4275), .ZN(n3267) );
  NAND4_X1 U4120 ( .A1(n3286), .A2(n3287), .A3(n3268), .A4(n3267), .ZN(n3270)
         );
  AOI21_X2 U4121 ( .B1(n3270), .B2(STATE2_REG_0__SCAN_IN), .A(n3269), .ZN(
        n3299) );
  NOR2_X1 U4122 ( .A1(n3999), .A2(n4465), .ZN(n3271) );
  NOR2_X1 U4123 ( .A1(n4047), .A2(n5190), .ZN(n3272) );
  AND2_X1 U4124 ( .A1(n4116), .A2(n4236), .ZN(n4056) );
  NAND2_X1 U4125 ( .A1(n4235), .A2(n4056), .ZN(n4066) );
  OAI211_X1 U4126 ( .C1(n3987), .C2(n3273), .A(n4066), .B(n4243), .ZN(n3274)
         );
  NAND2_X1 U4127 ( .A1(n3274), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3280) );
  INV_X1 U4128 ( .A(n4129), .ZN(n6499) );
  XNOR2_X1 U4129 ( .A(n4761), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5756)
         );
  NAND2_X1 U4130 ( .A1(n6499), .A2(n5756), .ZN(n3276) );
  INV_X1 U4131 ( .A(n3410), .ZN(n3303) );
  NAND2_X1 U4132 ( .A1(n3303), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3275) );
  AND2_X1 U4133 ( .A1(n3276), .A2(n3275), .ZN(n3277) );
  OAI211_X1 U4134 ( .C1(n3299), .C2(n5404), .A(n3280), .B(n3277), .ZN(n3297)
         );
  INV_X1 U4135 ( .A(n3277), .ZN(n3278) );
  NOR2_X1 U4136 ( .A1(n3278), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3279)
         );
  NAND2_X1 U4137 ( .A1(n3297), .A2(n2951), .ZN(n3377) );
  INV_X1 U4138 ( .A(n3377), .ZN(n3296) );
  INV_X1 U4139 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3281) );
  OR2_X2 U4140 ( .A1(n3299), .A2(n3281), .ZN(n3283) );
  MUX2_X1 U4141 ( .A(n3410), .B(n4129), .S(n4761), .Z(n3282) );
  NAND2_X1 U4142 ( .A1(n3283), .A2(n3282), .ZN(n3327) );
  INV_X1 U4143 ( .A(n3993), .ZN(n3285) );
  INV_X1 U4144 ( .A(n4247), .ZN(n3991) );
  NAND2_X1 U4145 ( .A1(n4116), .A2(n4065), .ZN(n3284) );
  AOI21_X1 U4146 ( .B1(n3285), .B2(n4006), .A(n4288), .ZN(n3294) );
  OR2_X1 U4147 ( .A1(n3286), .A2(n4000), .ZN(n4084) );
  INV_X1 U4148 ( .A(n3287), .ZN(n3292) );
  INV_X1 U4149 ( .A(n4001), .ZN(n3290) );
  NAND2_X1 U4150 ( .A1(n5900), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6408) );
  AOI21_X1 U4151 ( .B1(n4355), .B2(n3187), .A(n6408), .ZN(n3289) );
  NAND2_X1 U4152 ( .A1(n4247), .A2(n4697), .ZN(n3288) );
  OAI211_X1 U4153 ( .C1(n3290), .C2(n4236), .A(n3289), .B(n3288), .ZN(n3291)
         );
  NOR2_X1 U4154 ( .A1(n3292), .A2(n3291), .ZN(n3293) );
  OAI211_X1 U4155 ( .C1(n4284), .C2(n3294), .A(n4084), .B(n3293), .ZN(n3328)
         );
  INV_X1 U4156 ( .A(n3376), .ZN(n3295) );
  AND2_X2 U4157 ( .A1(n3298), .A2(n3297), .ZN(n3306) );
  INV_X1 U4158 ( .A(n3299), .ZN(n3408) );
  NAND2_X1 U4159 ( .A1(n3408), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3305) );
  AND2_X1 U4160 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3300) );
  NAND2_X1 U4161 ( .A1(n3300), .A2(n6376), .ZN(n6253) );
  INV_X1 U4162 ( .A(n3300), .ZN(n3301) );
  NAND2_X1 U4163 ( .A1(n3301), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3302) );
  NAND2_X1 U4164 ( .A1(n6253), .A2(n3302), .ZN(n4417) );
  AOI22_X1 U4165 ( .A1(n6499), .A2(n4417), .B1(n3303), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3304) );
  INV_X1 U4166 ( .A(n3306), .ZN(n3309) );
  INV_X1 U4167 ( .A(n3307), .ZN(n3308) );
  AOI22_X1 U4168 ( .A1(n3930), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3126), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4169 ( .A1(n3337), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3330), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4170 ( .A1(n3716), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4171 ( .A1(n3934), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3758), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3314) );
  NAND4_X1 U4172 ( .A1(n3317), .A2(n3316), .A3(n3315), .A4(n3314), .ZN(n3324)
         );
  BUF_X1 U4173 ( .A(n3318), .Z(n3914) );
  AOI22_X1 U4174 ( .A1(n3914), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3322) );
  INV_X1 U4175 ( .A(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n6584) );
  AOI22_X1 U4176 ( .A1(n3931), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3321) );
  AOI22_X1 U4177 ( .A1(n3942), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4178 ( .A1(n3944), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3319) );
  NAND4_X1 U4179 ( .A1(n3322), .A2(n3321), .A3(n3320), .A4(n3319), .ZN(n3323)
         );
  OAI22_X2 U4180 ( .A1(n4894), .A2(STATE2_REG_0__SCAN_IN), .B1(n4347), .B2(
        n4109), .ZN(n3326) );
  INV_X1 U4181 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5725) );
  OAI22_X1 U4182 ( .A1(n3501), .A2(n5725), .B1(n4347), .B2(n3361), .ZN(n3325)
         );
  CLKBUF_X1 U4183 ( .A(n3362), .Z(n3330) );
  AOI22_X1 U4184 ( .A1(n3330), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4186 ( .A1(n3331), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3126), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3335) );
  BUF_X1 U4187 ( .A(n3332), .Z(n3942) );
  AOI22_X1 U4188 ( .A1(n3930), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4189 ( .A1(n3914), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3333) );
  NAND4_X1 U4190 ( .A1(n3336), .A2(n3335), .A3(n3334), .A4(n3333), .ZN(n3345)
         );
  BUF_X1 U4191 ( .A(n3337), .Z(n3828) );
  AOI22_X1 U4192 ( .A1(n3716), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3828), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3343) );
  AOI22_X1 U4193 ( .A1(n3941), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3342) );
  BUF_X1 U4194 ( .A(n3338), .Z(n3758) );
  AOI22_X1 U4195 ( .A1(n3758), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3341) );
  BUF_X1 U4196 ( .A(n3339), .Z(n3931) );
  AOI22_X1 U4197 ( .A1(n3931), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3340) );
  NAND4_X1 U4198 ( .A1(n3343), .A2(n3342), .A3(n3341), .A4(n3340), .ZN(n3344)
         );
  INV_X1 U4199 ( .A(n4696), .ZN(n3360) );
  AOI22_X1 U4200 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3934), .B1(n3931), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3349) );
  AOI22_X1 U4201 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n3716), .B1(n3940), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3348) );
  AOI22_X1 U4202 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n3828), .B1(n3758), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3347) );
  AOI22_X1 U4203 ( .A1(n3836), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3346) );
  NAND4_X1 U4204 ( .A1(n3349), .A2(n3348), .A3(n3347), .A4(n3346), .ZN(n3355)
         );
  AOI22_X1 U4205 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n3330), .B1(n3941), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4206 ( .A1(n3823), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3352) );
  AOI22_X1 U4207 ( .A1(n3914), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3351) );
  AOI22_X1 U4208 ( .A1(n3930), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3350) );
  NAND4_X1 U4209 ( .A1(n3353), .A2(n3352), .A3(n3351), .A4(n3350), .ZN(n3354)
         );
  XNOR2_X1 U4210 ( .A(n3360), .B(n4354), .ZN(n3356) );
  NAND2_X1 U4211 ( .A1(n3356), .A2(n4239), .ZN(n3395) );
  INV_X1 U4212 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5717) );
  AOI21_X1 U4213 ( .B1(n4262), .B2(n4696), .A(n6520), .ZN(n3358) );
  NAND2_X1 U4214 ( .A1(n4299), .A2(n4354), .ZN(n3357) );
  OAI211_X1 U4215 ( .C1(n3501), .C2(n5717), .A(n3358), .B(n3357), .ZN(n3393)
         );
  NAND2_X1 U4216 ( .A1(n3394), .A2(n3393), .ZN(n3359) );
  NAND2_X1 U4217 ( .A1(n4239), .A2(n4696), .ZN(n4692) );
  INV_X1 U4218 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U4219 ( .A1(n4239), .A2(n3360), .ZN(n3375) );
  INV_X1 U4220 ( .A(n3361), .ZN(n3373) );
  AOI22_X1 U4221 ( .A1(n3934), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3828), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4222 ( .A1(n3330), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3365) );
  AOI22_X1 U4223 ( .A1(n3931), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4224 ( .A1(n3941), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3363) );
  NAND4_X1 U4225 ( .A1(n3366), .A2(n3365), .A3(n3364), .A4(n3363), .ZN(n3372)
         );
  AOI22_X1 U4226 ( .A1(n3930), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3126), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4227 ( .A1(n3716), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3758), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4228 ( .A1(n3914), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4229 ( .A1(n3942), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3367) );
  NAND4_X1 U4230 ( .A1(n3370), .A2(n3369), .A3(n3368), .A4(n3367), .ZN(n3371)
         );
  OR2_X1 U4231 ( .A1(n3372), .A2(n3371), .ZN(n4353) );
  NAND2_X1 U4232 ( .A1(n3373), .A2(n4353), .ZN(n3374) );
  OAI211_X1 U4233 ( .C1(n3501), .C2(n5721), .A(n3375), .B(n3374), .ZN(n3383)
         );
  XNOR2_X1 U4234 ( .A(n3377), .B(n3376), .ZN(n4886) );
  NAND2_X1 U4235 ( .A1(n4886), .A2(n6520), .ZN(n3379) );
  NAND2_X1 U4236 ( .A1(n4239), .A2(n4353), .ZN(n3378) );
  NAND2_X1 U4237 ( .A1(n3379), .A2(n3378), .ZN(n3386) );
  OAI21_X1 U4238 ( .B1(n3385), .B2(n3383), .A(n3386), .ZN(n3381) );
  NAND2_X1 U4239 ( .A1(n3385), .A2(n3383), .ZN(n3380) );
  NOR2_X2 U4240 ( .A1(n4236), .A2(n6405), .ZN(n3631) );
  NAND2_X1 U4241 ( .A1(n4346), .A2(n3631), .ZN(n3382) );
  NAND2_X1 U4242 ( .A1(n3382), .A2(n3885), .ZN(n3405) );
  INV_X1 U4243 ( .A(n3383), .ZN(n3384) );
  XNOR2_X1 U4244 ( .A(n3385), .B(n3384), .ZN(n3388) );
  INV_X1 U4245 ( .A(n3386), .ZN(n3387) );
  XNOR2_X1 U4246 ( .A(n3388), .B(n3387), .ZN(n4266) );
  NAND2_X1 U4247 ( .A1(n4266), .A2(n3631), .ZN(n3392) );
  AOI22_X1 U4248 ( .A1(n3669), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6405), .ZN(n3390) );
  AND2_X1 U4249 ( .A1(n4056), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3402) );
  NAND2_X1 U4250 ( .A1(n3402), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3389) );
  AND2_X1 U4251 ( .A1(n3390), .A2(n3389), .ZN(n3391) );
  NAND2_X1 U4252 ( .A1(n3392), .A2(n3391), .ZN(n4125) );
  AOI21_X1 U4253 ( .B1(n4615), .B2(n4292), .A(n6405), .ZN(n4119) );
  INV_X1 U4254 ( .A(n4654), .ZN(n6256) );
  NAND2_X1 U4255 ( .A1(n6256), .A2(n3631), .ZN(n3399) );
  AOI22_X1 U4256 ( .A1(n3669), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6405), .ZN(n3397) );
  NAND2_X1 U4257 ( .A1(n3402), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3396) );
  AND2_X1 U4258 ( .A1(n3397), .A2(n3396), .ZN(n3398) );
  NAND2_X1 U4259 ( .A1(n3399), .A2(n3398), .ZN(n4118) );
  NAND2_X1 U4260 ( .A1(n4119), .A2(n4118), .ZN(n4117) );
  INV_X1 U4261 ( .A(n4118), .ZN(n3400) );
  INV_X1 U4262 ( .A(n3650), .ZN(n3954) );
  INV_X1 U4263 ( .A(n3954), .ZN(n3961) );
  NAND2_X1 U4264 ( .A1(n3400), .A2(n3961), .ZN(n3401) );
  NAND2_X1 U4265 ( .A1(n4117), .A2(n3401), .ZN(n4126) );
  INV_X1 U4266 ( .A(n3402), .ZN(n3456) );
  OAI21_X1 U4267 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3441), .ZN(n6119) );
  AOI22_X1 U4268 ( .A1(n3668), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n3650), 
        .B2(n6119), .ZN(n3404) );
  NAND2_X1 U4269 ( .A1(n4238), .A2(EAX_REG_2__SCAN_IN), .ZN(n3403) );
  OAI211_X1 U4270 ( .C1(n3456), .C2(n5157), .A(n3404), .B(n3403), .ZN(n4148)
         );
  NAND2_X1 U4271 ( .A1(n4147), .A2(n4148), .ZN(n3407) );
  NAND2_X1 U4272 ( .A1(n3405), .A2(n4123), .ZN(n3406) );
  NAND2_X2 U4273 ( .A1(n3407), .A2(n3406), .ZN(n4153) );
  NAND2_X1 U4274 ( .A1(n3408), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3413) );
  NOR3_X1 U4275 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6376), .A3(n6372), 
        .ZN(n4612) );
  NAND2_X1 U4276 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4612), .ZN(n4517) );
  NAND2_X1 U4277 ( .A1(n6383), .A2(n4517), .ZN(n3409) );
  NAND3_X1 U4278 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4412) );
  INV_X1 U4279 ( .A(n4412), .ZN(n4272) );
  NAND2_X1 U4280 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4272), .ZN(n4306) );
  NAND2_X1 U4281 ( .A1(n3409), .A2(n4306), .ZN(n5755) );
  OAI22_X1 U4282 ( .A1(n4129), .A2(n5755), .B1(n3410), .B2(n6383), .ZN(n3411)
         );
  INV_X1 U4283 ( .A(n3411), .ZN(n3412) );
  INV_X1 U4284 ( .A(n3501), .ZN(n3424) );
  AOI22_X1 U4285 ( .A1(n3930), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3126), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3417) );
  AOI22_X1 U4286 ( .A1(n3828), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3330), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3416) );
  AOI22_X1 U4287 ( .A1(n3716), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3415) );
  AOI22_X1 U4288 ( .A1(n3934), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3758), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3414) );
  NAND4_X1 U4289 ( .A1(n3417), .A2(n3416), .A3(n3415), .A4(n3414), .ZN(n3423)
         );
  AOI22_X1 U4290 ( .A1(n3914), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3842), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3421) );
  AOI22_X1 U4291 ( .A1(n3931), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3420) );
  AOI22_X1 U4292 ( .A1(n3942), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3419) );
  AOI22_X1 U4293 ( .A1(n3944), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3418) );
  NAND4_X1 U4294 ( .A1(n3421), .A2(n3420), .A3(n3419), .A4(n3418), .ZN(n3422)
         );
  OR2_X1 U4295 ( .A1(n3423), .A2(n3422), .ZN(n4372) );
  AOI22_X1 U4296 ( .A1(n3424), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3499), 
        .B2(n4372), .ZN(n3425) );
  NAND2_X2 U4297 ( .A1(n3426), .A2(n3425), .ZN(n5696) );
  INV_X1 U4298 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5733) );
  OR2_X1 U4299 ( .A1(n3501), .A2(n5733), .ZN(n3440) );
  AOI22_X1 U4300 ( .A1(n3828), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3432) );
  BUF_X1 U4301 ( .A(n3126), .Z(n3836) );
  AOI22_X1 U4302 ( .A1(n3758), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4303 ( .A1(n3330), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4304 ( .A1(n3941), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3429) );
  NAND4_X1 U4305 ( .A1(n3432), .A2(n3431), .A3(n3430), .A4(n3429), .ZN(n3438)
         );
  AOI22_X1 U4306 ( .A1(n3716), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3930), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3436) );
  AOI22_X1 U4307 ( .A1(n3914), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3435) );
  AOI22_X1 U4308 ( .A1(n3934), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3434) );
  AOI22_X1 U4309 ( .A1(n3931), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3433) );
  NAND4_X1 U4310 ( .A1(n3436), .A2(n3435), .A3(n3434), .A4(n3433), .ZN(n3437)
         );
  OR2_X1 U4311 ( .A1(n3438), .A2(n3437), .ZN(n4389) );
  NAND2_X1 U4312 ( .A1(n3499), .A2(n4389), .ZN(n3439) );
  NAND2_X1 U4313 ( .A1(n3440), .A2(n3439), .ZN(n3475) );
  XNOR2_X1 U4314 ( .A(n3496), .B(n3475), .ZN(n4371) );
  AOI21_X1 U4315 ( .B1(n4663), .B2(n3452), .A(n3471), .ZN(n4667) );
  NAND2_X1 U4316 ( .A1(n6405), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3443)
         );
  NAND2_X1 U4317 ( .A1(n4238), .A2(EAX_REG_4__SCAN_IN), .ZN(n3442) );
  OAI211_X1 U4318 ( .C1(n3456), .C2(n6607), .A(n3443), .B(n3442), .ZN(n3444)
         );
  NAND2_X1 U4319 ( .A1(n3444), .A2(n3954), .ZN(n3445) );
  OAI21_X1 U4320 ( .B1(n4667), .B2(n3954), .A(n3445), .ZN(n3446) );
  AOI21_X1 U4321 ( .B1(n4371), .B2(n3631), .A(n3446), .ZN(n4140) );
  INV_X1 U4322 ( .A(n3447), .ZN(n3449) );
  NAND2_X1 U4323 ( .A1(n3449), .A2(n3448), .ZN(n3450) );
  NAND2_X1 U4324 ( .A1(n3450), .A2(n4486), .ZN(n3451) );
  AND2_X2 U4325 ( .A1(n3451), .A2(n3496), .ZN(n4832) );
  OAI21_X1 U4326 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3453), .A(n3452), 
        .ZN(n6108) );
  AOI22_X1 U4327 ( .A1(n3961), .A2(n6108), .B1(n3668), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3455) );
  NAND2_X1 U4328 ( .A1(n4238), .A2(EAX_REG_3__SCAN_IN), .ZN(n3454) );
  OAI211_X1 U4329 ( .C1(n3456), .C2(n4206), .A(n3455), .B(n3454), .ZN(n3457)
         );
  NAND2_X1 U4331 ( .A1(n3476), .A2(n3475), .ZN(n3470) );
  INV_X1 U4332 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5737) );
  AOI22_X1 U4333 ( .A1(n3930), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3462) );
  AOI22_X1 U4334 ( .A1(n3828), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3330), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3461) );
  AOI22_X1 U4335 ( .A1(n3716), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3460) );
  AOI22_X1 U4336 ( .A1(n3934), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3758), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3459) );
  NAND4_X1 U4337 ( .A1(n3462), .A2(n3461), .A3(n3460), .A4(n3459), .ZN(n3468)
         );
  AOI22_X1 U4338 ( .A1(n3914), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3941), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4339 ( .A1(n3931), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3465) );
  AOI22_X1 U4340 ( .A1(n3942), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4341 ( .A1(n3944), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3463) );
  NAND4_X1 U4342 ( .A1(n3466), .A2(n3465), .A3(n3464), .A4(n3463), .ZN(n3467)
         );
  OR2_X1 U4343 ( .A1(n3468), .A2(n3467), .ZN(n4390) );
  NAND2_X1 U4344 ( .A1(n3499), .A2(n4390), .ZN(n3469) );
  OAI21_X1 U4345 ( .B1(n3501), .B2(n5737), .A(n3469), .ZN(n3474) );
  XNOR2_X1 U4346 ( .A(n3470), .B(n3474), .ZN(n4379) );
  INV_X1 U4347 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4309) );
  OAI21_X1 U4348 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3471), .A(n3504), 
        .ZN(n6100) );
  AOI22_X1 U4349 ( .A1(n3650), .A2(n6100), .B1(n3668), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3472) );
  OAI21_X1 U4350 ( .B1(n3956), .B2(n4309), .A(n3472), .ZN(n3473) );
  AND2_X1 U4351 ( .A1(n3475), .A2(n3474), .ZN(n3498) );
  NAND2_X1 U4352 ( .A1(n3476), .A2(n3498), .ZN(n3490) );
  INV_X1 U4353 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5741) );
  OR2_X1 U4354 ( .A1(n3501), .A2(n5741), .ZN(n3488) );
  AOI22_X1 U4355 ( .A1(n3930), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3480) );
  AOI22_X1 U4356 ( .A1(n3828), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3330), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4357 ( .A1(n3716), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4358 ( .A1(n3934), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3758), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3477) );
  NAND4_X1 U4359 ( .A1(n3480), .A2(n3479), .A3(n3478), .A4(n3477), .ZN(n3486)
         );
  AOI22_X1 U4360 ( .A1(n3914), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3842), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3484) );
  AOI22_X1 U4361 ( .A1(n3931), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4362 ( .A1(n3332), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4363 ( .A1(n3944), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3481) );
  NAND4_X1 U4364 ( .A1(n3484), .A2(n3483), .A3(n3482), .A4(n3481), .ZN(n3485)
         );
  OR2_X1 U4365 ( .A1(n3486), .A2(n3485), .ZN(n4679) );
  NAND2_X1 U4366 ( .A1(n3499), .A2(n4679), .ZN(n3487) );
  NAND2_X1 U4367 ( .A1(n3488), .A2(n3487), .ZN(n3497) );
  INV_X1 U4368 ( .A(n3497), .ZN(n3489) );
  NAND2_X1 U4369 ( .A1(n4238), .A2(EAX_REG_6__SCAN_IN), .ZN(n3492) );
  INV_X1 U4370 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6305) );
  OAI21_X1 U4371 ( .B1(n6305), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6405), 
        .ZN(n3491) );
  XNOR2_X1 U4372 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n3504), .ZN(n4475) );
  AOI22_X1 U4373 ( .A1(n3492), .A2(n3491), .B1(n3650), .B2(n4475), .ZN(n3493)
         );
  INV_X1 U4374 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5749) );
  NAND2_X1 U4375 ( .A1(n3499), .A2(n4696), .ZN(n3500) );
  OAI21_X1 U4376 ( .B1(n3501), .B2(n5749), .A(n3500), .ZN(n3502) );
  INV_X1 U4377 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3509) );
  INV_X1 U4378 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3503) );
  OR2_X1 U4379 ( .A1(n3505), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3506) );
  NAND2_X1 U4380 ( .A1(n3506), .A2(n3525), .ZN(n6092) );
  NAND2_X1 U4381 ( .A1(n6092), .A2(n3961), .ZN(n3508) );
  NAND2_X1 U4382 ( .A1(n3669), .A2(EAX_REG_7__SCAN_IN), .ZN(n3507) );
  OAI211_X1 U4383 ( .C1(n3509), .C2(n3885), .A(n3508), .B(n3507), .ZN(n3510)
         );
  NOR2_X2 U4384 ( .A1(n4595), .A2(n4594), .ZN(n4582) );
  INV_X1 U4385 ( .A(n3631), .ZN(n3673) );
  AOI22_X1 U4386 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3828), .B1(n3931), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4387 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n3940), .B1(n3330), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4388 ( .A1(n3914), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4389 ( .A1(n3758), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3511) );
  NAND4_X1 U4390 ( .A1(n3514), .A2(n3513), .A3(n3512), .A4(n3511), .ZN(n3520)
         );
  AOI22_X1 U4391 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n3934), .B1(n3842), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3518) );
  AOI22_X1 U4392 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n3716), .B1(n3836), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4393 ( .A1(n3942), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3516) );
  AOI22_X1 U4394 ( .A1(n3930), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3515) );
  NAND4_X1 U4395 ( .A1(n3518), .A2(n3517), .A3(n3516), .A4(n3515), .ZN(n3519)
         );
  NOR2_X1 U4396 ( .A1(n3520), .A2(n3519), .ZN(n3524) );
  XNOR2_X1 U4397 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3525), .ZN(n4713) );
  INV_X1 U4398 ( .A(n4713), .ZN(n3521) );
  AOI22_X1 U4399 ( .A1(n3668), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n3650), 
        .B2(n3521), .ZN(n3523) );
  NAND2_X1 U4400 ( .A1(n4238), .A2(EAX_REG_8__SCAN_IN), .ZN(n3522) );
  OAI211_X1 U4401 ( .C1(n3673), .C2(n3524), .A(n3523), .B(n3522), .ZN(n4581)
         );
  INV_X1 U4402 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3527) );
  XNOR2_X1 U4403 ( .A(n3542), .B(n3527), .ZN(n4919) );
  AOI22_X1 U4404 ( .A1(n3716), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3828), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3531) );
  AOI22_X1 U4405 ( .A1(n3934), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3530) );
  AOI22_X1 U4406 ( .A1(n3914), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U4407 ( .A1(n3942), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3528) );
  NAND4_X1 U4408 ( .A1(n3531), .A2(n3530), .A3(n3529), .A4(n3528), .ZN(n3537)
         );
  AOI22_X1 U4409 ( .A1(n3330), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3535) );
  AOI22_X1 U4410 ( .A1(n3930), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3758), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3534) );
  AOI22_X1 U4411 ( .A1(n3339), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4412 ( .A1(n3915), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3532) );
  NAND4_X1 U4413 ( .A1(n3535), .A2(n3534), .A3(n3533), .A4(n3532), .ZN(n3536)
         );
  OAI21_X1 U4414 ( .B1(n3537), .B2(n3536), .A(n3631), .ZN(n3540) );
  NAND2_X1 U4415 ( .A1(n4238), .A2(EAX_REG_9__SCAN_IN), .ZN(n3539) );
  NAND2_X1 U4416 ( .A1(n3668), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3538)
         );
  NAND3_X1 U4417 ( .A1(n3540), .A2(n3539), .A3(n3538), .ZN(n3541) );
  AOI21_X1 U4418 ( .B1(n4919), .B2(n3650), .A(n3541), .ZN(n4720) );
  XOR2_X1 U4419 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3558), .Z(n5957) );
  INV_X1 U4420 ( .A(n5957), .ZN(n4955) );
  AOI22_X1 U4421 ( .A1(n3934), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3914), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3546) );
  AOI22_X1 U4422 ( .A1(n3330), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3545) );
  AOI22_X1 U4423 ( .A1(n3823), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4424 ( .A1(n3915), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3543) );
  NAND4_X1 U4425 ( .A1(n3546), .A2(n3545), .A3(n3544), .A4(n3543), .ZN(n3552)
         );
  AOI22_X1 U4426 ( .A1(n3828), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3930), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4427 ( .A1(n3716), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4428 ( .A1(n3758), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4429 ( .A1(n3931), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3547) );
  NAND4_X1 U4430 ( .A1(n3550), .A2(n3549), .A3(n3548), .A4(n3547), .ZN(n3551)
         );
  OAI21_X1 U4431 ( .B1(n3552), .B2(n3551), .A(n3631), .ZN(n3555) );
  NAND2_X1 U4432 ( .A1(n4238), .A2(EAX_REG_10__SCAN_IN), .ZN(n3554) );
  NAND2_X1 U4433 ( .A1(n3668), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3553)
         );
  NAND3_X1 U4434 ( .A1(n3555), .A2(n3554), .A3(n3553), .ZN(n3556) );
  AOI21_X1 U4435 ( .B1(n4955), .B2(n3650), .A(n3556), .ZN(n4920) );
  NAND2_X1 U4436 ( .A1(n3558), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3574)
         );
  INV_X1 U4437 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3559) );
  XNOR2_X1 U4438 ( .A(n3574), .B(n3559), .ZN(n5008) );
  AOI22_X1 U4439 ( .A1(n3339), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3842), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4440 ( .A1(n3331), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4441 ( .A1(n3930), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4442 ( .A1(n3318), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3560) );
  NAND4_X1 U4443 ( .A1(n3563), .A2(n3562), .A3(n3561), .A4(n3560), .ZN(n3569)
         );
  AOI22_X1 U4444 ( .A1(n3716), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3330), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3567) );
  AOI22_X1 U4445 ( .A1(n3828), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3758), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4446 ( .A1(n3944), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4447 ( .A1(n3942), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3564) );
  NAND4_X1 U4448 ( .A1(n3567), .A2(n3566), .A3(n3565), .A4(n3564), .ZN(n3568)
         );
  OAI21_X1 U4449 ( .B1(n3569), .B2(n3568), .A(n3631), .ZN(n3572) );
  NAND2_X1 U4450 ( .A1(n4238), .A2(EAX_REG_11__SCAN_IN), .ZN(n3571) );
  NAND2_X1 U4451 ( .A1(n3668), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3570)
         );
  NAND3_X1 U4452 ( .A1(n3572), .A2(n3571), .A3(n3570), .ZN(n3573) );
  AOI21_X1 U4453 ( .B1(n5008), .B2(n3961), .A(n3573), .ZN(n4982) );
  XOR2_X1 U4454 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3588), .Z(n5133) );
  AOI22_X1 U4455 ( .A1(n3914), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3578) );
  AOI22_X1 U4456 ( .A1(n3716), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3330), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3577) );
  AOI22_X1 U4457 ( .A1(n3930), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4458 ( .A1(n3828), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3575) );
  NAND4_X1 U4459 ( .A1(n3578), .A2(n3577), .A3(n3576), .A4(n3575), .ZN(n3584)
         );
  AOI22_X1 U4460 ( .A1(n3934), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4461 ( .A1(n3758), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4462 ( .A1(n3915), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3732), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4463 ( .A1(n3823), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3579) );
  NAND4_X1 U4464 ( .A1(n3582), .A2(n3581), .A3(n3580), .A4(n3579), .ZN(n3583)
         );
  OR2_X1 U4465 ( .A1(n3584), .A2(n3583), .ZN(n3585) );
  AOI22_X1 U4466 ( .A1(n3631), .A2(n3585), .B1(n3668), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3587) );
  NAND2_X1 U4467 ( .A1(n3669), .A2(EAX_REG_12__SCAN_IN), .ZN(n3586) );
  OAI211_X1 U4468 ( .C1(n5133), .C2(n3954), .A(n3587), .B(n3586), .ZN(n5014)
         );
  NAND2_X1 U4469 ( .A1(n3588), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3589)
         );
  INV_X1 U4470 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6533) );
  NAND2_X1 U4471 ( .A1(n3589), .A2(n6533), .ZN(n3590) );
  NAND2_X1 U4472 ( .A1(n3590), .A2(n3607), .ZN(n5947) );
  NAND2_X1 U4473 ( .A1(n5947), .A2(n3961), .ZN(n3593) );
  NOR2_X1 U4474 ( .A1(n3885), .A2(n6533), .ZN(n3591) );
  AOI21_X1 U4475 ( .B1(n4238), .B2(EAX_REG_13__SCAN_IN), .A(n3591), .ZN(n3592)
         );
  NAND2_X1 U4476 ( .A1(n3593), .A2(n3592), .ZN(n3605) );
  XNOR2_X2 U4477 ( .A(n5013), .B(n3605), .ZN(n5119) );
  AOI22_X1 U4478 ( .A1(n3331), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3716), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4479 ( .A1(n3339), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4480 ( .A1(n3362), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4481 ( .A1(n3914), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3594) );
  NAND4_X1 U4482 ( .A1(n3597), .A2(n3596), .A3(n3595), .A4(n3594), .ZN(n3603)
         );
  AOI22_X1 U4483 ( .A1(n3915), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4484 ( .A1(n3828), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4485 ( .A1(n3930), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3599) );
  AOI22_X1 U4486 ( .A1(n3338), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3598) );
  NAND4_X1 U4487 ( .A1(n3601), .A2(n3600), .A3(n3599), .A4(n3598), .ZN(n3602)
         );
  OR2_X1 U4488 ( .A1(n3603), .A2(n3602), .ZN(n3604) );
  AND2_X1 U4489 ( .A1(n3631), .A2(n3604), .ZN(n5118) );
  INV_X1 U4490 ( .A(n3605), .ZN(n3606) );
  INV_X1 U4491 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6566) );
  NAND2_X1 U4492 ( .A1(n3665), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3648)
         );
  INV_X1 U4493 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5166) );
  INV_X1 U4494 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3608) );
  XNOR2_X1 U4495 ( .A(n3694), .B(n3608), .ZN(n5586) );
  AOI22_X1 U4496 ( .A1(n4238), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6405), .ZN(n3622) );
  AOI22_X1 U4497 ( .A1(n3716), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3930), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4498 ( .A1(n3931), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4499 ( .A1(n3915), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4500 ( .A1(n3914), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3609) );
  NAND4_X1 U4501 ( .A1(n3612), .A2(n3611), .A3(n3610), .A4(n3609), .ZN(n3620)
         );
  AOI22_X1 U4502 ( .A1(n3330), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3338), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4503 ( .A1(n3934), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3732), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4504 ( .A1(n3828), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3616) );
  NAND2_X1 U4505 ( .A1(n3940), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3614) );
  AOI21_X1 U4506 ( .B1(n3822), .B2(INSTQUEUE_REG_9__2__SCAN_IN), .A(n3961), 
        .ZN(n3613) );
  AND2_X1 U4507 ( .A1(n3614), .A2(n3613), .ZN(n3615) );
  NAND4_X1 U4508 ( .A1(n3618), .A2(n3617), .A3(n3616), .A4(n3615), .ZN(n3619)
         );
  NOR2_X1 U4509 ( .A1(n4006), .A2(n6520), .ZN(n3958) );
  NAND2_X1 U4510 ( .A1(n3924), .A2(n3954), .ZN(n3768) );
  OAI21_X1 U4511 ( .B1(n3620), .B2(n3619), .A(n3768), .ZN(n3621) );
  AOI22_X1 U4512 ( .A1(n5586), .A2(n3961), .B1(n3622), .B2(n3621), .ZN(n5453)
         );
  AOI22_X1 U4513 ( .A1(n3362), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4514 ( .A1(n3914), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3732), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4515 ( .A1(n3339), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4516 ( .A1(n3331), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3623) );
  NAND4_X1 U4517 ( .A1(n3626), .A2(n3625), .A3(n3624), .A4(n3623), .ZN(n3633)
         );
  AOI22_X1 U4518 ( .A1(n3828), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3842), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4519 ( .A1(n3716), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4520 ( .A1(n3758), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4521 ( .A1(n3930), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3627) );
  NAND4_X1 U4522 ( .A1(n3630), .A2(n3629), .A3(n3628), .A4(n3627), .ZN(n3632)
         );
  OAI21_X1 U4523 ( .B1(n3633), .B2(n3632), .A(n3631), .ZN(n3637) );
  NAND2_X1 U4524 ( .A1(n3669), .A2(EAX_REG_15__SCAN_IN), .ZN(n3636) );
  XOR2_X1 U4525 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3665), .Z(n5592) );
  INV_X1 U4526 ( .A(n5592), .ZN(n3634) );
  AOI22_X1 U4527 ( .A1(n3668), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n3650), 
        .B2(n3634), .ZN(n3635) );
  AND3_X1 U4528 ( .A1(n3637), .A2(n3636), .A3(n3635), .ZN(n5173) );
  AOI22_X1 U4529 ( .A1(n3914), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3330), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4530 ( .A1(n3716), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4531 ( .A1(n3428), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4532 ( .A1(n3930), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3638) );
  NAND4_X1 U4533 ( .A1(n3641), .A2(n3640), .A3(n3639), .A4(n3638), .ZN(n3647)
         );
  AOI22_X1 U4534 ( .A1(n3931), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4535 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n3828), .B1(n3758), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4536 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n3934), .B1(n3942), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4537 ( .A1(n3915), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3732), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3642) );
  NAND4_X1 U4538 ( .A1(n3645), .A2(n3644), .A3(n3643), .A4(n3642), .ZN(n3646)
         );
  OR2_X1 U4539 ( .A1(n3647), .A2(n3646), .ZN(n3654) );
  INV_X1 U4540 ( .A(EAX_REG_16__SCAN_IN), .ZN(n3652) );
  INV_X1 U4541 ( .A(n3648), .ZN(n3649) );
  XNOR2_X1 U4542 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3649), .ZN(n5244)
         );
  AOI22_X1 U4543 ( .A1(n3650), .A2(n5244), .B1(n3668), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3651) );
  OAI21_X1 U4544 ( .B1(n3956), .B2(n3652), .A(n3651), .ZN(n3653) );
  AOI21_X1 U4545 ( .B1(n3958), .B2(n3654), .A(n3653), .ZN(n5148) );
  NOR2_X1 U4546 ( .A1(n5173), .A2(n5148), .ZN(n3674) );
  AOI22_X1 U4547 ( .A1(n3931), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4548 ( .A1(n3828), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3330), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4549 ( .A1(n3942), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3732), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4550 ( .A1(n3338), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3655) );
  NAND4_X1 U4551 ( .A1(n3658), .A2(n3657), .A3(n3656), .A4(n3655), .ZN(n3664)
         );
  AOI22_X1 U4552 ( .A1(n3934), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3842), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4553 ( .A1(n3716), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U4554 ( .A1(n3318), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4555 ( .A1(n3930), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3659) );
  NAND4_X1 U4556 ( .A1(n3662), .A2(n3661), .A3(n3660), .A4(n3659), .ZN(n3663)
         );
  NOR2_X1 U4557 ( .A1(n3664), .A2(n3663), .ZN(n3672) );
  INV_X1 U4558 ( .A(n3665), .ZN(n3666) );
  OAI21_X1 U4559 ( .B1(PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n3667), .A(n3666), 
        .ZN(n5603) );
  AOI22_X1 U4560 ( .A1(n3961), .A2(n5603), .B1(n3668), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3671) );
  NAND2_X1 U4561 ( .A1(n3669), .A2(EAX_REG_14__SCAN_IN), .ZN(n3670) );
  OAI211_X1 U4562 ( .C1(n3673), .C2(n3672), .A(n3671), .B(n3670), .ZN(n5474)
         );
  AND2_X1 U4563 ( .A1(n3674), .A2(n5474), .ZN(n5149) );
  INV_X1 U4564 ( .A(n3694), .ZN(n3677) );
  OR2_X1 U4565 ( .A1(n3675), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3676)
         );
  NAND2_X1 U4566 ( .A1(n3677), .A2(n3676), .ZN(n5937) );
  AOI22_X1 U4567 ( .A1(n3828), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3930), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4568 ( .A1(n3716), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3330), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4569 ( .A1(n3338), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3679) );
  AOI22_X1 U4570 ( .A1(n3318), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3732), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3678) );
  NAND4_X1 U4571 ( .A1(n3681), .A2(n3680), .A3(n3679), .A4(n3678), .ZN(n3687)
         );
  AOI22_X1 U4572 ( .A1(n3931), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3842), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4573 ( .A1(n3940), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4574 ( .A1(n3331), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4575 ( .A1(n3428), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3682) );
  NAND4_X1 U4576 ( .A1(n3685), .A2(n3684), .A3(n3683), .A4(n3682), .ZN(n3686)
         );
  NOR2_X1 U4577 ( .A1(n3687), .A2(n3686), .ZN(n3688) );
  NOR2_X1 U4578 ( .A1(n3924), .A2(n3688), .ZN(n3692) );
  INV_X1 U4579 ( .A(EAX_REG_17__SCAN_IN), .ZN(n3690) );
  NAND2_X1 U4580 ( .A1(n6405), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3689)
         );
  OAI211_X1 U4581 ( .C1(n3956), .C2(n3690), .A(n3954), .B(n3689), .ZN(n3691)
         );
  OAI22_X1 U4582 ( .A1(n5937), .A2(n3954), .B1(n3692), .B2(n3691), .ZN(n5521)
         );
  INV_X1 U4583 ( .A(n5521), .ZN(n3693) );
  AND2_X1 U4584 ( .A1(n5149), .A2(n3693), .ZN(n5450) );
  INV_X1 U4585 ( .A(n5451), .ZN(n3712) );
  OR2_X1 U4586 ( .A1(n3695), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3696)
         );
  NAND2_X1 U4587 ( .A1(n3696), .A2(n3747), .ZN(n5861) );
  AOI22_X1 U4588 ( .A1(n3931), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3915), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4589 ( .A1(n3331), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3828), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4590 ( .A1(n3318), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3698) );
  AOI22_X1 U4591 ( .A1(n3940), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3697) );
  NAND4_X1 U4592 ( .A1(n3700), .A2(n3699), .A3(n3698), .A4(n3697), .ZN(n3706)
         );
  AOI22_X1 U4593 ( .A1(n3716), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3758), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4594 ( .A1(n3362), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4595 ( .A1(n3930), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3732), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4596 ( .A1(n3823), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3701) );
  NAND4_X1 U4597 ( .A1(n3704), .A2(n3703), .A3(n3702), .A4(n3701), .ZN(n3705)
         );
  NOR2_X1 U4598 ( .A1(n3706), .A2(n3705), .ZN(n3707) );
  NOR2_X1 U4599 ( .A1(n3924), .A2(n3707), .ZN(n3711) );
  INV_X1 U4600 ( .A(EAX_REG_19__SCAN_IN), .ZN(n3709) );
  NAND2_X1 U4601 ( .A1(n6405), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3708)
         );
  OAI211_X1 U4602 ( .C1(n3956), .C2(n3709), .A(n3954), .B(n3708), .ZN(n3710)
         );
  OAI22_X1 U4603 ( .A1(n5861), .A2(n3954), .B1(n3711), .B2(n3710), .ZN(n5516)
         );
  NOR2_X1 U4604 ( .A1(n3712), .A2(n5516), .ZN(n5176) );
  INV_X1 U4605 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5445) );
  INV_X1 U4606 ( .A(n3770), .ZN(n3715) );
  OR2_X1 U4607 ( .A1(n3713), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3714)
         );
  NAND2_X1 U4608 ( .A1(n3715), .A2(n3714), .ZN(n5852) );
  OR2_X1 U4609 ( .A1(n5852), .A2(n3954), .ZN(n3731) );
  AOI22_X1 U4610 ( .A1(n3934), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3914), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4611 ( .A1(n3716), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3330), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4612 ( .A1(n3828), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3758), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4613 ( .A1(n3944), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3717) );
  NAND4_X1 U4614 ( .A1(n3720), .A2(n3719), .A3(n3718), .A4(n3717), .ZN(n3726)
         );
  AOI22_X1 U4615 ( .A1(n3931), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3915), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4616 ( .A1(n3940), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4617 ( .A1(n3930), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4618 ( .A1(n3428), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3721) );
  NAND4_X1 U4619 ( .A1(n3724), .A2(n3723), .A3(n3722), .A4(n3721), .ZN(n3725)
         );
  NOR2_X1 U4620 ( .A1(n3726), .A2(n3725), .ZN(n3729) );
  OAI21_X1 U4621 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6305), .A(n6405), 
        .ZN(n3728) );
  NAND2_X1 U4622 ( .A1(n4238), .A2(EAX_REG_21__SCAN_IN), .ZN(n3727) );
  OAI211_X1 U4623 ( .C1(n3924), .C2(n3729), .A(n3728), .B(n3727), .ZN(n3730)
         );
  NAND2_X1 U4624 ( .A1(n3731), .A2(n3730), .ZN(n5504) );
  INV_X1 U4625 ( .A(n5504), .ZN(n3750) );
  AOI22_X1 U4626 ( .A1(n3930), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4627 ( .A1(n3915), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3338), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4628 ( .A1(n3332), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3732), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4629 ( .A1(n3828), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3733) );
  NAND4_X1 U4630 ( .A1(n3736), .A2(n3735), .A3(n3734), .A4(n3733), .ZN(n3744)
         );
  AOI22_X1 U4631 ( .A1(n3914), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4632 ( .A1(n3940), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4633 ( .A1(n3934), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3740) );
  NAND2_X1 U4634 ( .A1(n3716), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3738)
         );
  AOI21_X1 U4635 ( .B1(n3822), .B2(INSTQUEUE_REG_9__4__SCAN_IN), .A(n3961), 
        .ZN(n3737) );
  AND2_X1 U4636 ( .A1(n3738), .A2(n3737), .ZN(n3739) );
  NAND4_X1 U4637 ( .A1(n3742), .A2(n3741), .A3(n3740), .A4(n3739), .ZN(n3743)
         );
  OAI21_X1 U4638 ( .B1(n3744), .B2(n3743), .A(n3768), .ZN(n3746) );
  AOI22_X1 U4639 ( .A1(n4238), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6405), .ZN(n3745) );
  NAND2_X1 U4640 ( .A1(n3746), .A2(n3745), .ZN(n3749) );
  XNOR2_X1 U4641 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n3747), .ZN(n5565)
         );
  NAND2_X1 U4642 ( .A1(n3961), .A2(n5565), .ZN(n3748) );
  NAND2_X1 U4643 ( .A1(n3749), .A2(n3748), .ZN(n5441) );
  INV_X1 U4644 ( .A(n5441), .ZN(n5501) );
  AND2_X1 U4645 ( .A1(n3750), .A2(n5501), .ZN(n5175) );
  INV_X1 U4646 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5303) );
  XNOR2_X1 U4647 ( .A(n3770), .B(n5303), .ZN(n5307) );
  AOI22_X1 U4648 ( .A1(n3940), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4649 ( .A1(n3331), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4650 ( .A1(n3915), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3755) );
  NAND2_X1 U4651 ( .A1(n3716), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3753)
         );
  AOI21_X1 U4652 ( .B1(n3822), .B2(INSTQUEUE_REG_9__6__SCAN_IN), .A(n3961), 
        .ZN(n3752) );
  AND2_X1 U4653 ( .A1(n3753), .A2(n3752), .ZN(n3754) );
  NAND4_X1 U4654 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3764)
         );
  AOI22_X1 U4655 ( .A1(n3930), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4656 ( .A1(n3318), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3758), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4657 ( .A1(n3931), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4658 ( .A1(n3828), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3759) );
  NAND4_X1 U4659 ( .A1(n3762), .A2(n3761), .A3(n3760), .A4(n3759), .ZN(n3763)
         );
  OR2_X1 U4660 ( .A1(n3764), .A2(n3763), .ZN(n3767) );
  INV_X1 U4661 ( .A(EAX_REG_22__SCAN_IN), .ZN(n3765) );
  OAI22_X1 U4662 ( .A1(n3956), .A2(n3765), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5303), .ZN(n3766) );
  AOI21_X1 U4663 ( .B1(n3768), .B2(n3767), .A(n3766), .ZN(n3769) );
  AOI21_X1 U4664 ( .B1(n5307), .B2(n3961), .A(n3769), .ZN(n5213) );
  INV_X1 U4665 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5274) );
  NAND2_X1 U4666 ( .A1(n3881), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3871)
         );
  INV_X1 U4667 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5312) );
  INV_X1 U4668 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3852) );
  XNOR2_X1 U4669 ( .A(n3902), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5199)
         );
  INV_X1 U4670 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5181) );
  NOR2_X1 U4671 ( .A1(n5181), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3771) );
  AOI211_X1 U4672 ( .C1(n4238), .C2(EAX_REG_28__SCAN_IN), .A(n3961), .B(n3771), 
        .ZN(n3851) );
  AOI22_X1 U4673 ( .A1(n3930), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3126), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4674 ( .A1(n3337), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4675 ( .A1(n3716), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4676 ( .A1(n3331), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3338), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3772) );
  NAND4_X1 U4677 ( .A1(n3775), .A2(n3774), .A3(n3773), .A4(n3772), .ZN(n3781)
         );
  AOI22_X1 U4678 ( .A1(n3318), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3842), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4679 ( .A1(n3931), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3935), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4680 ( .A1(n3332), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4681 ( .A1(n3944), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3776) );
  NAND4_X1 U4682 ( .A1(n3779), .A2(n3778), .A3(n3777), .A4(n3776), .ZN(n3780)
         );
  OR2_X1 U4683 ( .A1(n3781), .A2(n3780), .ZN(n3907) );
  AOI22_X1 U4684 ( .A1(n3318), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3915), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4685 ( .A1(n3934), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3126), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4686 ( .A1(n3337), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3758), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4687 ( .A1(n3931), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3782) );
  NAND4_X1 U4688 ( .A1(n3785), .A2(n3784), .A3(n3783), .A4(n3782), .ZN(n3791)
         );
  AOI22_X1 U4689 ( .A1(n3930), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4690 ( .A1(n3716), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4691 ( .A1(n3428), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3935), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4692 ( .A1(n3332), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3786) );
  NAND4_X1 U4693 ( .A1(n3789), .A2(n3788), .A3(n3787), .A4(n3786), .ZN(n3790)
         );
  NOR2_X1 U4694 ( .A1(n3791), .A2(n3790), .ZN(n3855) );
  AOI22_X1 U4695 ( .A1(n3915), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4696 ( .A1(n3716), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4697 ( .A1(n3330), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3758), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4698 ( .A1(n3914), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3792) );
  NAND4_X1 U4699 ( .A1(n3795), .A2(n3794), .A3(n3793), .A4(n3792), .ZN(n3801)
         );
  AOI22_X1 U4700 ( .A1(n3934), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3828), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4701 ( .A1(n3823), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3935), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4702 ( .A1(n3931), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4703 ( .A1(n3930), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3796) );
  NAND4_X1 U4704 ( .A1(n3799), .A2(n3798), .A3(n3797), .A4(n3796), .ZN(n3800)
         );
  NOR2_X1 U4705 ( .A1(n3801), .A2(n3800), .ZN(n3883) );
  AOI22_X1 U4706 ( .A1(n3930), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3842), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4707 ( .A1(n3716), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3330), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4708 ( .A1(n3934), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4709 ( .A1(n3332), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3802) );
  NAND4_X1 U4710 ( .A1(n3805), .A2(n3804), .A3(n3803), .A4(n3802), .ZN(n3811)
         );
  AOI22_X1 U4711 ( .A1(n3337), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4712 ( .A1(n3914), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4713 ( .A1(n3758), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4714 ( .A1(n3931), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3935), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3806) );
  NAND4_X1 U4715 ( .A1(n3809), .A2(n3808), .A3(n3807), .A4(n3806), .ZN(n3810)
         );
  NOR2_X1 U4716 ( .A1(n3811), .A2(n3810), .ZN(n3872) );
  AOI22_X1 U4717 ( .A1(n3931), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3930), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4718 ( .A1(n3716), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4719 ( .A1(n3337), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3758), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4720 ( .A1(n3332), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3935), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3812) );
  NAND4_X1 U4721 ( .A1(n3815), .A2(n3814), .A3(n3813), .A4(n3812), .ZN(n3821)
         );
  AOI22_X1 U4722 ( .A1(n3934), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3330), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4723 ( .A1(n3915), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4724 ( .A1(n3944), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4725 ( .A1(n3914), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3816) );
  NAND4_X1 U4726 ( .A1(n3819), .A2(n3818), .A3(n3817), .A4(n3816), .ZN(n3820)
         );
  NOR2_X1 U4727 ( .A1(n3821), .A2(n3820), .ZN(n3892) );
  AOI22_X1 U4728 ( .A1(n3931), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3915), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4729 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n3934), .B1(n3914), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4730 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3330), .B1(n3758), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4731 ( .A1(n3823), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3824) );
  NAND4_X1 U4732 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3835)
         );
  AOI22_X1 U4733 ( .A1(n3716), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4734 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n3828), .B1(n3836), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4735 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n3930), .B1(n3942), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4736 ( .A1(n3944), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3830) );
  NAND4_X1 U4737 ( .A1(n3833), .A2(n3832), .A3(n3831), .A4(n3830), .ZN(n3834)
         );
  NOR2_X1 U4738 ( .A1(n3835), .A2(n3834), .ZN(n3893) );
  OR2_X1 U4739 ( .A1(n3892), .A2(n3893), .ZN(n3884) );
  NOR3_X1 U4740 ( .A1(n3883), .A2(n3872), .A3(n3884), .ZN(n3864) );
  AOI22_X1 U4741 ( .A1(n3930), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4742 ( .A1(n3337), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3330), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4743 ( .A1(n3716), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4744 ( .A1(n3934), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3758), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3838) );
  NAND4_X1 U4745 ( .A1(n3841), .A2(n3840), .A3(n3839), .A4(n3838), .ZN(n3848)
         );
  AOI22_X1 U4746 ( .A1(n3914), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3842), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4747 ( .A1(n3339), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3935), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4748 ( .A1(n3332), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4749 ( .A1(n3944), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3843) );
  NAND4_X1 U4750 ( .A1(n3846), .A2(n3845), .A3(n3844), .A4(n3843), .ZN(n3847)
         );
  OR2_X1 U4751 ( .A1(n3848), .A2(n3847), .ZN(n3862) );
  NAND2_X1 U4752 ( .A1(n3864), .A2(n3862), .ZN(n3856) );
  NOR2_X1 U4753 ( .A1(n3855), .A2(n3856), .ZN(n3908) );
  XOR2_X1 U4754 ( .A(n3907), .B(n3908), .Z(n3849) );
  NAND2_X1 U4755 ( .A1(n3849), .A2(n3958), .ZN(n3850) );
  AOI22_X1 U4756 ( .A1(n5199), .A2(n3961), .B1(n3851), .B2(n3850), .ZN(n5180)
         );
  NAND2_X1 U4757 ( .A1(n3853), .A2(n3852), .ZN(n3854) );
  NAND2_X1 U4758 ( .A1(n3902), .A2(n3854), .ZN(n5813) );
  XNOR2_X1 U4759 ( .A(n3856), .B(n3855), .ZN(n3857) );
  NOR2_X1 U4760 ( .A1(n3857), .A2(n3924), .ZN(n3861) );
  INV_X1 U4761 ( .A(EAX_REG_27__SCAN_IN), .ZN(n3859) );
  NAND2_X1 U4762 ( .A1(n6405), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3858)
         );
  OAI211_X1 U4763 ( .C1(n3956), .C2(n3859), .A(n3954), .B(n3858), .ZN(n3860)
         );
  OAI22_X1 U4764 ( .A1(n5813), .A2(n3954), .B1(n3861), .B2(n3860), .ZN(n5206)
         );
  XNOR2_X1 U4765 ( .A(n3871), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5330)
         );
  INV_X1 U4766 ( .A(n3862), .ZN(n3863) );
  XNOR2_X1 U4767 ( .A(n3864), .B(n3863), .ZN(n3868) );
  INV_X1 U4768 ( .A(EAX_REG_26__SCAN_IN), .ZN(n3866) );
  NAND2_X1 U4769 ( .A1(n6405), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3865)
         );
  OAI211_X1 U4770 ( .C1(n3956), .C2(n3866), .A(n3954), .B(n3865), .ZN(n3867)
         );
  AOI21_X1 U4771 ( .B1(n3868), .B2(n3958), .A(n3867), .ZN(n3869) );
  AOI21_X1 U4772 ( .B1(n5330), .B2(n3961), .A(n3869), .ZN(n5316) );
  INV_X1 U4773 ( .A(n5316), .ZN(n3900) );
  OR2_X1 U4774 ( .A1(n3881), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3870)
         );
  AND2_X1 U4775 ( .A1(n3871), .A2(n3870), .ZN(n5826) );
  NAND2_X1 U4776 ( .A1(n5826), .A2(n3961), .ZN(n3880) );
  NOR2_X1 U4777 ( .A1(n3884), .A2(n3883), .ZN(n3873) );
  XNOR2_X1 U4778 ( .A(n3873), .B(n3872), .ZN(n3874) );
  NAND2_X1 U4779 ( .A1(n3874), .A2(n3958), .ZN(n3878) );
  NAND2_X1 U4780 ( .A1(n6405), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3875)
         );
  NAND2_X1 U4781 ( .A1(n3954), .A2(n3875), .ZN(n3876) );
  AOI21_X1 U4782 ( .B1(n4238), .B2(EAX_REG_25__SCAN_IN), .A(n3876), .ZN(n3877)
         );
  NAND2_X1 U4783 ( .A1(n3878), .A2(n3877), .ZN(n3879) );
  NAND2_X1 U4784 ( .A1(n3880), .A2(n3879), .ZN(n5283) );
  AND2_X1 U4785 ( .A1(n3890), .A2(n5274), .ZN(n3882) );
  OR2_X1 U4786 ( .A1(n3882), .A2(n3881), .ZN(n5348) );
  XNOR2_X1 U4787 ( .A(n3884), .B(n3883), .ZN(n3888) );
  NOR2_X1 U4788 ( .A1(n3885), .A2(n5274), .ZN(n3886) );
  AOI21_X1 U4789 ( .B1(n4238), .B2(EAX_REG_24__SCAN_IN), .A(n3886), .ZN(n3887)
         );
  OAI21_X1 U4790 ( .B1(n3888), .B2(n3924), .A(n3887), .ZN(n3889) );
  AOI21_X1 U4791 ( .B1(n5348), .B2(n3961), .A(n3889), .ZN(n5267) );
  OAI21_X1 U4792 ( .B1(n3891), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n3890), 
        .ZN(n5844) );
  OR2_X1 U4793 ( .A1(n5844), .A2(n3954), .ZN(n3899) );
  XNOR2_X1 U4794 ( .A(n3893), .B(n3892), .ZN(n3897) );
  NAND2_X1 U4795 ( .A1(n6405), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3894)
         );
  NAND2_X1 U4796 ( .A1(n3954), .A2(n3894), .ZN(n3895) );
  AOI21_X1 U4797 ( .B1(n4238), .B2(EAX_REG_23__SCAN_IN), .A(n3895), .ZN(n3896)
         );
  OAI21_X1 U4798 ( .B1(n3924), .B2(n3897), .A(n3896), .ZN(n3898) );
  NAND2_X1 U4799 ( .A1(n3899), .A2(n3898), .ZN(n5257) );
  OR2_X1 U4800 ( .A1(n5267), .A2(n5257), .ZN(n5263) );
  OR2_X1 U4801 ( .A1(n5283), .A2(n5263), .ZN(n5280) );
  OR2_X1 U4802 ( .A1(n3900), .A2(n5280), .ZN(n5205) );
  NOR2_X1 U4803 ( .A1(n5206), .A2(n5205), .ZN(n5178) );
  AND2_X1 U4804 ( .A1(n5180), .A2(n5178), .ZN(n3901) );
  AND2_X1 U4805 ( .A1(n5213), .A2(n3901), .ZN(n5179) );
  NAND2_X1 U4806 ( .A1(n3903), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3965)
         );
  INV_X1 U4807 ( .A(n3903), .ZN(n3905) );
  INV_X1 U4808 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3904) );
  NAND2_X1 U4809 ( .A1(n3905), .A2(n3904), .ZN(n3906) );
  NAND2_X1 U4810 ( .A1(n3965), .A2(n3906), .ZN(n5554) );
  NAND2_X1 U4811 ( .A1(n3908), .A2(n3907), .ZN(n3928) );
  AOI22_X1 U4812 ( .A1(n3330), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4813 ( .A1(n3930), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3126), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4814 ( .A1(n3339), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4815 ( .A1(n3332), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3910) );
  NAND4_X1 U4816 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3921)
         );
  AOI22_X1 U4817 ( .A1(n3716), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3337), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4818 ( .A1(n3331), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3338), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4819 ( .A1(n3914), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3935), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4820 ( .A1(n3915), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3916) );
  NAND4_X1 U4821 ( .A1(n3919), .A2(n3918), .A3(n3917), .A4(n3916), .ZN(n3920)
         );
  NOR2_X1 U4822 ( .A1(n3921), .A2(n3920), .ZN(n3929) );
  XNOR2_X1 U4823 ( .A(n3928), .B(n3929), .ZN(n3925) );
  AOI21_X1 U4824 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6405), .A(n3961), 
        .ZN(n3923) );
  NAND2_X1 U4825 ( .A1(n4238), .A2(EAX_REG_29__SCAN_IN), .ZN(n3922) );
  OAI211_X1 U4826 ( .C1(n3925), .C2(n3924), .A(n3923), .B(n3922), .ZN(n3926)
         );
  OAI21_X1 U4827 ( .B1(n5554), .B2(n3954), .A(n3926), .ZN(n5428) );
  INV_X1 U4828 ( .A(n5428), .ZN(n3927) );
  AND2_X1 U4829 ( .A1(n5179), .A2(n3927), .ZN(n5375) );
  XNOR2_X1 U4830 ( .A(n3965), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5387)
         );
  NOR2_X1 U4831 ( .A1(n3929), .A2(n3928), .ZN(n3952) );
  AOI22_X1 U4832 ( .A1(n3931), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3930), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4833 ( .A1(n3716), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3337), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3938) );
  AOI22_X1 U4834 ( .A1(n3934), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3126), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4835 ( .A1(n3428), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3935), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3936) );
  NAND4_X1 U4836 ( .A1(n3939), .A2(n3938), .A3(n3937), .A4(n3936), .ZN(n3950)
         );
  AOI22_X1 U4837 ( .A1(n3362), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3940), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4838 ( .A1(n3941), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3338), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4839 ( .A1(n3318), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3942), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4840 ( .A1(n3944), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3943), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3945) );
  NAND4_X1 U4841 ( .A1(n3948), .A2(n3947), .A3(n3946), .A4(n3945), .ZN(n3949)
         );
  NOR2_X1 U4842 ( .A1(n3950), .A2(n3949), .ZN(n3951) );
  XNOR2_X1 U4843 ( .A(n3952), .B(n3951), .ZN(n3959) );
  INV_X1 U4844 ( .A(EAX_REG_30__SCAN_IN), .ZN(n3955) );
  NAND2_X1 U4845 ( .A1(n6405), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3953)
         );
  OAI211_X1 U4846 ( .C1(n3956), .C2(n3955), .A(n3954), .B(n3953), .ZN(n3957)
         );
  AOI21_X1 U4847 ( .B1(n3959), .B2(n3958), .A(n3957), .ZN(n3960) );
  AOI21_X1 U4848 ( .B1(n5387), .B2(n3961), .A(n3960), .ZN(n5376) );
  AND2_X1 U4849 ( .A1(n5375), .A2(n5376), .ZN(n3962) );
  NAND2_X1 U4850 ( .A1(n5502), .A2(n3962), .ZN(n3963) );
  XOR2_X1 U4851 ( .A(n3964), .B(n3963), .Z(n5423) );
  INV_X1 U4852 ( .A(n5423), .ZN(n3983) );
  INV_X1 U4853 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5379) );
  INV_X1 U4854 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3966) );
  XNOR2_X1 U4855 ( .A(n3967), .B(n3966), .ZN(n5418) );
  NAND2_X1 U4856 ( .A1(n4992), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4462) );
  NAND2_X1 U4857 ( .A1(n4284), .A2(n6422), .ZN(n4055) );
  AND3_X1 U4858 ( .A1(n4055), .A2(n3968), .A3(n3187), .ZN(n3969) );
  NAND3_X1 U4859 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n3972) );
  INV_X1 U4860 ( .A(REIP_REG_11__SCAN_IN), .ZN(n5017) );
  INV_X1 U4861 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6436) );
  NAND3_X1 U4862 ( .A1(REIP_REG_3__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n4605) );
  NOR2_X1 U4863 ( .A1(n6436), .A2(n4605), .ZN(n5979) );
  NAND2_X1 U4864 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5979), .ZN(n4456) );
  NAND2_X1 U4865 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n5967) );
  NOR2_X1 U4866 ( .A1(n4456), .A2(n5967), .ZN(n4585) );
  NAND2_X1 U4867 ( .A1(REIP_REG_8__SCAN_IN), .A2(n4585), .ZN(n4914) );
  NAND2_X1 U4868 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n4990) );
  NOR3_X1 U4869 ( .A1(n5017), .A2(n4914), .A3(n4990), .ZN(n4993) );
  NAND4_X1 U4870 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .A4(n4993), .ZN(n5469) );
  NOR2_X1 U4871 ( .A1(n5978), .A2(n5469), .ZN(n5160) );
  NAND4_X1 U4872 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_17__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .A4(n5160), .ZN(n5853) );
  NOR2_X1 U4873 ( .A1(n3972), .A2(n5853), .ZN(n5836) );
  NAND4_X1 U4874 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5836), .ZN(n5325) );
  INV_X1 U4875 ( .A(n5325), .ZN(n3971) );
  NAND3_X1 U4876 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n3975) );
  INV_X1 U4877 ( .A(n3975), .ZN(n3970) );
  NAND2_X1 U4878 ( .A1(n3971), .A2(n3970), .ZN(n5814) );
  NAND2_X1 U4879 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n3977) );
  NOR2_X1 U4880 ( .A1(n5384), .A2(REIP_REG_29__SCAN_IN), .ZN(n5437) );
  NOR2_X1 U4881 ( .A1(n4890), .A2(n5469), .ZN(n5161) );
  NAND4_X1 U4882 ( .A1(n5161), .A2(REIP_REG_15__SCAN_IN), .A3(
        REIP_REG_17__SCAN_IN), .A4(REIP_REG_16__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U4883 ( .A1(n5978), .A2(n4992), .ZN(n5459) );
  OAI21_X1 U4884 ( .B1(n5458), .B2(n3972), .A(n5459), .ZN(n5847) );
  INV_X1 U4885 ( .A(REIP_REG_22__SCAN_IN), .ZN(n5225) );
  INV_X1 U4886 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6457) );
  NOR2_X1 U4887 ( .A1(n5225), .A2(n6457), .ZN(n5837) );
  NAND2_X1 U4888 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5837), .ZN(n3973) );
  NAND2_X1 U4889 ( .A1(n5459), .A2(n3973), .ZN(n3974) );
  AND2_X1 U4890 ( .A1(n5847), .A2(n3974), .ZN(n5839) );
  NAND2_X1 U4891 ( .A1(n5459), .A2(n3975), .ZN(n3976) );
  AND2_X1 U4892 ( .A1(n5839), .A2(n3976), .ZN(n5816) );
  INV_X1 U4893 ( .A(n3977), .ZN(n3978) );
  OR2_X1 U4894 ( .A1(n5978), .A2(n3978), .ZN(n3979) );
  NAND2_X1 U4895 ( .A1(n5816), .A2(n3979), .ZN(n5439) );
  NOR2_X1 U4896 ( .A1(n5437), .A2(n5439), .ZN(n5390) );
  OAI21_X1 U4897 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5978), .A(n5390), .ZN(n3981) );
  INV_X1 U4898 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6473) );
  INV_X1 U4899 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6470) );
  NOR4_X1 U4900 ( .A1(n5384), .A2(REIP_REG_31__SCAN_IN), .A3(n6473), .A4(n6470), .ZN(n3980) );
  INV_X1 U4901 ( .A(n4697), .ZN(n6506) );
  NAND2_X1 U4902 ( .A1(n4299), .A2(n4047), .ZN(n4600) );
  NAND2_X1 U4903 ( .A1(n6506), .A2(n4600), .ZN(n3989) );
  NAND2_X1 U4904 ( .A1(n6483), .A2(n6405), .ZN(n6308) );
  OR2_X1 U4905 ( .A1(n6308), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5812) );
  INV_X1 U4906 ( .A(n5812), .ZN(n4470) );
  OAI21_X1 U4907 ( .B1(n4470), .B2(READREQUEST_REG_SCAN_IN), .A(n6503), .ZN(
        n3986) );
  OAI21_X1 U4908 ( .B1(n6503), .B2(n3989), .A(n3986), .ZN(U3474) );
  INV_X1 U4909 ( .A(n4026), .ZN(n4045) );
  OR2_X1 U4910 ( .A1(n4048), .A2(n4045), .ZN(n3988) );
  INV_X1 U4911 ( .A(n4107), .ZN(n4087) );
  NOR2_X1 U4912 ( .A1(n4047), .A2(n3187), .ZN(n4009) );
  INV_X1 U4913 ( .A(n4009), .ZN(n4599) );
  AOI22_X1 U4914 ( .A1(n3988), .A2(n3987), .B1(n4087), .B2(n4599), .ZN(n5906)
         );
  NAND2_X1 U4915 ( .A1(n3989), .A2(n6422), .ZN(n3990) );
  NAND2_X1 U4916 ( .A1(n3990), .A2(n6592), .ZN(n6504) );
  NAND2_X1 U4917 ( .A1(n5906), .A2(n6504), .ZN(n6389) );
  AND2_X1 U4918 ( .A1(n6389), .A2(n4053), .ZN(n5914) );
  INV_X1 U4919 ( .A(MORE_REG_SCAN_IN), .ZN(n4018) );
  AOI21_X1 U4920 ( .B1(n3991), .B2(n3187), .A(n4697), .ZN(n3992) );
  OR2_X1 U4921 ( .A1(n3993), .A2(n3992), .ZN(n4043) );
  AOI21_X1 U4922 ( .B1(n4056), .B2(n4299), .A(n4280), .ZN(n3994) );
  AOI21_X1 U4923 ( .B1(n3995), .B2(n5432), .A(n3994), .ZN(n3997) );
  NOR2_X1 U4924 ( .A1(n4600), .A2(n4049), .ZN(n4088) );
  OAI21_X1 U4925 ( .B1(n4088), .B2(n4068), .A(n4355), .ZN(n3996) );
  AND2_X1 U4926 ( .A1(n3997), .A2(n3996), .ZN(n3998) );
  AND2_X1 U4927 ( .A1(n4043), .A2(n3998), .ZN(n4086) );
  AND2_X1 U4928 ( .A1(n4299), .A2(n3999), .ZN(n4348) );
  INV_X1 U4929 ( .A(n4348), .ZN(n4038) );
  INV_X1 U4930 ( .A(n4000), .ZN(n4003) );
  NAND2_X1 U4931 ( .A1(n4235), .A2(n4292), .ZN(n4002) );
  INV_X1 U4932 ( .A(n4006), .ZN(n5394) );
  NAND2_X1 U4933 ( .A1(n5394), .A2(n4001), .ZN(n4210) );
  OAI211_X1 U4934 ( .C1(n4038), .C2(n4003), .A(n4002), .B(n4210), .ZN(n4004)
         );
  INV_X1 U4935 ( .A(n4004), .ZN(n4005) );
  AND3_X1 U4936 ( .A1(n4086), .A2(n4005), .A3(n4084), .ZN(n4072) );
  NOR2_X1 U4937 ( .A1(n4006), .A2(n4284), .ZN(n4042) );
  AND2_X1 U4938 ( .A1(n4006), .A2(n4299), .ZN(n4007) );
  NOR2_X1 U4939 ( .A1(n4011), .A2(n4007), .ZN(n4044) );
  AND2_X1 U4940 ( .A1(n4044), .A2(n4008), .ZN(n4127) );
  NAND2_X1 U4941 ( .A1(n5394), .A2(n4009), .ZN(n4010) );
  NOR2_X1 U4942 ( .A1(n4011), .A2(n4010), .ZN(n4232) );
  NOR3_X1 U4943 ( .A1(n4012), .A2(n4127), .A3(n4232), .ZN(n4014) );
  INV_X1 U4944 ( .A(n4048), .ZN(n4013) );
  OAI22_X1 U4945 ( .A1(n4014), .A2(n4107), .B1(n4045), .B2(n4013), .ZN(n4015)
         );
  AOI21_X1 U4946 ( .B1(n4196), .B2(n4107), .A(n4015), .ZN(n6388) );
  INV_X1 U4947 ( .A(n6388), .ZN(n4016) );
  NAND2_X1 U4948 ( .A1(n4016), .A2(n5914), .ZN(n4017) );
  OAI21_X1 U4949 ( .B1(n5914), .B2(n4018), .A(n4017), .ZN(U3471) );
  OR2_X1 U4950 ( .A1(n4091), .A2(n6506), .ZN(n6398) );
  INV_X1 U4951 ( .A(n6398), .ZN(n4019) );
  NAND2_X1 U4952 ( .A1(n4020), .A2(n6075), .ZN(n6082) );
  AOI22_X1 U4953 ( .A1(n6073), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6079), .ZN(n4021) );
  INV_X1 U4954 ( .A(DATAI_5_), .ZN(n4276) );
  OR2_X1 U4955 ( .A1(n6058), .A2(n4276), .ZN(n4166) );
  NAND2_X1 U4956 ( .A1(n4021), .A2(n4166), .ZN(U2929) );
  AOI22_X1 U4957 ( .A1(n6073), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6079), .ZN(n4022) );
  INV_X1 U4958 ( .A(n6058), .ZN(n6080) );
  NAND2_X1 U4959 ( .A1(n6080), .A2(DATAI_3_), .ZN(n4170) );
  NAND2_X1 U4960 ( .A1(n4022), .A2(n4170), .ZN(U2927) );
  AOI22_X1 U4961 ( .A1(n6073), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6079), .ZN(n4023) );
  NAND2_X1 U4962 ( .A1(n6080), .A2(DATAI_2_), .ZN(n4173) );
  NAND2_X1 U4963 ( .A1(n4023), .A2(n4173), .ZN(U2926) );
  AOI22_X1 U4964 ( .A1(n6073), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n6079), .ZN(n4024) );
  NAND2_X1 U4965 ( .A1(n6080), .A2(DATAI_1_), .ZN(n4161) );
  NAND2_X1 U4966 ( .A1(n4024), .A2(n4161), .ZN(U2925) );
  AOI22_X1 U4967 ( .A1(n6073), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6079), .ZN(n4025) );
  NAND2_X1 U4968 ( .A1(n6080), .A2(DATAI_4_), .ZN(n4164) );
  NAND2_X1 U4969 ( .A1(n4025), .A2(n4164), .ZN(U2928) );
  INV_X1 U4970 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6050) );
  AND2_X1 U4971 ( .A1(n4026), .A2(n4047), .ZN(n6366) );
  NAND2_X1 U4972 ( .A1(n4233), .A2(n6366), .ZN(n4027) );
  NAND2_X1 U4973 ( .A1(n6075), .A2(n4027), .ZN(n4029) );
  NAND2_X1 U4974 ( .A1(n6020), .A2(n3187), .ZN(n4195) );
  NAND2_X1 U4975 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4228) );
  NOR2_X1 U4976 ( .A1(n4228), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6041) );
  INV_X1 U4977 ( .A(n6041), .ZN(n6395) );
  INV_X1 U4978 ( .A(n6395), .ZN(n6501) );
  AOI22_X1 U4979 ( .A1(n6501), .A2(UWORD_REG_9__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4030) );
  OAI21_X1 U4980 ( .B1(n6050), .B2(n4195), .A(n4030), .ZN(U2898) );
  AOI22_X1 U4981 ( .A1(n6501), .A2(UWORD_REG_10__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4031) );
  OAI21_X1 U4982 ( .B1(n3866), .B2(n4195), .A(n4031), .ZN(U2897) );
  INV_X1 U4983 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6047) );
  AOI22_X1 U4984 ( .A1(n6501), .A2(UWORD_REG_8__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4032) );
  OAI21_X1 U4985 ( .B1(n6047), .B2(n4195), .A(n4032), .ZN(U2899) );
  INV_X1 U4986 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6609) );
  AOI22_X1 U4987 ( .A1(n6501), .A2(UWORD_REG_12__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4033) );
  OAI21_X1 U4988 ( .B1(n6609), .B2(n4195), .A(n4033), .ZN(U2895) );
  INV_X1 U4989 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U4990 ( .A1(n6501), .A2(UWORD_REG_13__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4034) );
  OAI21_X1 U4991 ( .B1(n4035), .B2(n4195), .A(n4034), .ZN(U2894) );
  AOI22_X1 U4992 ( .A1(n6501), .A2(UWORD_REG_11__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4036) );
  OAI21_X1 U4993 ( .B1(n3859), .B2(n4195), .A(n4036), .ZN(U2896) );
  AOI22_X1 U4994 ( .A1(n6501), .A2(UWORD_REG_14__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4037) );
  OAI21_X1 U4995 ( .B1(n3955), .B2(n4195), .A(n4037), .ZN(U2893) );
  INV_X2 U4996 ( .A(n4615), .ZN(n4766) );
  INV_X1 U4997 ( .A(n4691), .ZN(n4676) );
  NAND2_X1 U4998 ( .A1(n4766), .A2(n4676), .ZN(n4041) );
  OAI21_X1 U4999 ( .B1(n6506), .B2(n4354), .A(n4038), .ZN(n4039) );
  INV_X1 U5000 ( .A(n4039), .ZN(n4040) );
  NAND2_X1 U5001 ( .A1(n4041), .A2(n4040), .ZN(n4362) );
  XNOR2_X1 U5002 ( .A(n4362), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4139)
         );
  INV_X1 U5003 ( .A(n4042), .ZN(n4052) );
  NAND2_X1 U5004 ( .A1(n4044), .A2(n4043), .ZN(n4046) );
  NAND2_X1 U5005 ( .A1(n4046), .A2(n4045), .ZN(n4090) );
  NAND2_X1 U5006 ( .A1(n4047), .A2(n6422), .ZN(n4050) );
  NOR2_X1 U5007 ( .A1(READY_N), .A2(n4048), .ZN(n4094) );
  NAND3_X1 U5008 ( .A1(n4050), .A2(n4094), .A3(n4049), .ZN(n4051) );
  OAI211_X1 U5009 ( .C1(n4052), .C2(n4107), .A(n4090), .B(n4051), .ZN(n4054)
         );
  NAND2_X1 U5010 ( .A1(n4054), .A2(n4053), .ZN(n4060) );
  INV_X1 U5011 ( .A(READY_N), .ZN(n6592) );
  NAND2_X1 U5012 ( .A1(n4055), .A2(n6592), .ZN(n4057) );
  INV_X1 U5013 ( .A(n4056), .ZN(n5192) );
  OAI211_X1 U5014 ( .C1(n4091), .C2(n4057), .A(n3187), .B(n5192), .ZN(n4058)
         );
  NAND3_X1 U5015 ( .A1(n4233), .A2(n4058), .A3(n4280), .ZN(n4059) );
  INV_X1 U5016 ( .A(n4127), .ZN(n6387) );
  NOR2_X1 U5017 ( .A1(n4066), .A2(n4262), .ZN(n4061) );
  NOR2_X1 U5018 ( .A1(n4232), .A2(n4061), .ZN(n4063) );
  OR2_X1 U5019 ( .A1(n4091), .A2(n4092), .ZN(n4062) );
  NAND4_X1 U5020 ( .A1(n6387), .A2(n4063), .A3(n4243), .A4(n4062), .ZN(n4064)
         );
  OAI21_X1 U5021 ( .B1(n4066), .B2(n4065), .A(n6398), .ZN(n4067) );
  AND2_X2 U5022 ( .A1(n4077), .A2(n4067), .ZN(n6168) );
  NOR2_X1 U5023 ( .A1(n4068), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4069)
         );
  OR2_X1 U5024 ( .A1(n4070), .A2(n4069), .ZN(n4653) );
  INV_X1 U5025 ( .A(n4653), .ZN(n4071) );
  INV_X1 U5026 ( .A(n5585), .ZN(n6167) );
  AND2_X1 U5027 ( .A1(n6167), .A2(REIP_REG_0__SCAN_IN), .ZN(n4136) );
  AOI21_X1 U5028 ( .B1(n6168), .B2(n4071), .A(n4136), .ZN(n4080) );
  INV_X1 U5029 ( .A(n4072), .ZN(n4073) );
  AND2_X1 U5030 ( .A1(n4077), .A2(n4073), .ZN(n4823) );
  INV_X1 U5031 ( .A(n4823), .ZN(n4074) );
  OR2_X1 U5032 ( .A1(n4967), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4076)
         );
  OR2_X1 U5033 ( .A1(n4077), .A2(n6167), .ZN(n4075) );
  NAND2_X1 U5034 ( .A1(n4076), .A2(n4075), .ZN(n5685) );
  INV_X1 U5035 ( .A(n4967), .ZN(n4078) );
  OAI22_X1 U5036 ( .A1(n5685), .A2(n4965), .B1(n4078), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4079) );
  OAI211_X1 U5037 ( .C1(n4139), .C2(n5680), .A(n4080), .B(n4079), .ZN(U3018)
         );
  INV_X1 U5038 ( .A(n4081), .ZN(n4082) );
  NOR2_X1 U5039 ( .A1(n4082), .A2(n4235), .ZN(n4083) );
  AND2_X1 U5040 ( .A1(n4091), .A2(n4083), .ZN(n4085) );
  AND4_X1 U5041 ( .A1(n4086), .A2(n4085), .A3(n4243), .A4(n4084), .ZN(n5397)
         );
  INV_X1 U5042 ( .A(n5397), .ZN(n4205) );
  AOI22_X1 U5043 ( .A1(n6256), .A2(n4205), .B1(n5394), .B2(n6369), .ZN(n6367)
         );
  INV_X1 U5044 ( .A(n5900), .ZN(n6486) );
  NOR2_X1 U5045 ( .A1(n6367), .A2(n6486), .ZN(n4104) );
  INV_X1 U5046 ( .A(n5399), .ZN(n6484) );
  NAND2_X1 U5047 ( .A1(n4196), .A2(n4087), .ZN(n4100) );
  INV_X1 U5048 ( .A(n4088), .ZN(n4089) );
  AND2_X1 U5049 ( .A1(n4090), .A2(n4089), .ZN(n4098) );
  AOI21_X1 U5050 ( .B1(n4092), .B2(n6422), .A(READY_N), .ZN(n4093) );
  OAI211_X1 U5051 ( .C1(n6366), .C2(n3188), .A(n4093), .B(n4107), .ZN(n4097)
         );
  NAND2_X1 U5052 ( .A1(n4232), .A2(n4107), .ZN(n4096) );
  INV_X1 U5053 ( .A(n4094), .ZN(n4234) );
  OR2_X1 U5054 ( .A1(n4243), .A2(n4234), .ZN(n4095) );
  AND4_X1 U5055 ( .A1(n4098), .A2(n4097), .A3(n4096), .A4(n4095), .ZN(n4099)
         );
  OR2_X1 U5056 ( .A1(n6520), .A2(n4228), .ZN(n6480) );
  INV_X1 U5057 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5913) );
  OAI22_X1 U5058 ( .A1(n6375), .A2(n6407), .B1(n6480), .B2(n5913), .ZN(n5899)
         );
  NAND2_X1 U5059 ( .A1(n6520), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6481) );
  INV_X1 U5060 ( .A(n6481), .ZN(n4101) );
  NOR2_X1 U5061 ( .A1(n5899), .A2(n4101), .ZN(n6488) );
  INV_X1 U5062 ( .A(n6488), .ZN(n5904) );
  OAI21_X1 U5063 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6484), .A(n5904), 
        .ZN(n4102) );
  INV_X1 U5064 ( .A(n4102), .ZN(n5403) );
  OAI21_X1 U5065 ( .B1(n4237), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n5403), 
        .ZN(n4103) );
  OAI22_X1 U5066 ( .A1(n4104), .A2(n4103), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5904), .ZN(n4106) );
  NAND3_X1 U5067 ( .A1(n6366), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n5900), .ZN(n4105) );
  NAND2_X1 U5068 ( .A1(n4106), .A2(n4105), .ZN(U3461) );
  NOR2_X1 U5069 ( .A1(n4107), .A2(n6407), .ZN(n4108) );
  NAND2_X1 U5070 ( .A1(n4196), .A2(n4108), .ZN(n4115) );
  NAND2_X1 U5071 ( .A1(n4288), .A2(n4236), .ZN(n4110) );
  NOR2_X1 U5072 ( .A1(n4110), .A2(n4109), .ZN(n4113) );
  NOR2_X1 U5073 ( .A1(n5190), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4111) );
  AND2_X1 U5074 ( .A1(n4111), .A2(n4280), .ZN(n4112) );
  NAND4_X1 U5075 ( .A1(n4113), .A2(n4121), .A3(n4238), .A4(n4112), .ZN(n4114)
         );
  INV_X1 U5076 ( .A(n4116), .ZN(n5422) );
  NAND2_X2 U5077 ( .A1(n5532), .A2(n5422), .ZN(n5535) );
  OAI21_X1 U5078 ( .B1(n4119), .B2(n4118), .A(n4117), .ZN(n4659) );
  OAI222_X1 U5079 ( .A1(n4653), .A2(n5535), .B1(n5532), .B2(n4120), .C1(n2945), 
        .C2(n4659), .ZN(U2859) );
  XNOR2_X1 U5080 ( .A(n4122), .B(n4121), .ZN(n5682) );
  INV_X1 U5081 ( .A(n4123), .ZN(n4124) );
  OAI21_X1 U5082 ( .B1(n4126), .B2(n4125), .A(n4124), .ZN(n4889) );
  OAI222_X1 U5083 ( .A1(n5682), .A2(n5535), .B1(n5532), .B2(n3010), .C1(n2945), 
        .C2(n4889), .ZN(U2858) );
  INV_X1 U5084 ( .A(n4659), .ZN(n4137) );
  NAND3_X1 U5085 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), 
        .A3(n6520), .ZN(n6415) );
  INV_X1 U5086 ( .A(n6415), .ZN(n4128) );
  NAND2_X1 U5087 ( .A1(n6500), .A2(n4128), .ZN(n5591) );
  NAND2_X1 U5088 ( .A1(n4129), .A2(n6308), .ZN(n4130) );
  NAND2_X1 U5089 ( .A1(n4130), .A2(n6520), .ZN(n4131) );
  INV_X1 U5090 ( .A(n6109), .ZN(n5597) );
  NAND2_X1 U5091 ( .A1(n6520), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4133) );
  NAND2_X1 U5092 ( .A1(n6305), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4132) );
  AND2_X1 U5093 ( .A1(n4133), .A2(n4132), .ZN(n4407) );
  INV_X1 U5094 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4134) );
  AOI21_X1 U5095 ( .B1(n5597), .B2(n4407), .A(n4134), .ZN(n4135) );
  AOI211_X1 U5096 ( .C1(n4137), .C2(n2946), .A(n4136), .B(n4135), .ZN(n4138)
         );
  OAI21_X1 U5097 ( .B1(n4139), .B2(n5912), .A(n4138), .ZN(U2986) );
  INV_X1 U5098 ( .A(n4153), .ZN(n4146) );
  OAI21_X1 U5099 ( .B1(n4146), .B2(n4152), .A(n4140), .ZN(n4141) );
  NAND2_X1 U5100 ( .A1(n4141), .A2(n4259), .ZN(n4664) );
  OR2_X1 U5101 ( .A1(n4142), .A2(n4154), .ZN(n4143) );
  NAND2_X1 U5102 ( .A1(n4143), .A2(n4254), .ZN(n4603) );
  OAI22_X1 U5103 ( .A1(n5535), .A2(n4603), .B1(n6594), .B2(n5532), .ZN(n4144)
         );
  INV_X1 U5104 ( .A(n4144), .ZN(n4145) );
  OAI21_X1 U5105 ( .B1(n4664), .B2(n2945), .A(n4145), .ZN(U2855) );
  OAI21_X1 U5106 ( .B1(n4148), .B2(n4147), .A(n4146), .ZN(n6110) );
  XOR2_X1 U5107 ( .A(n4150), .B(n4149), .Z(n6169) );
  INV_X1 U5108 ( .A(n5535), .ZN(n5511) );
  AOI22_X1 U5109 ( .A1(n6169), .A2(n5511), .B1(n5509), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4151) );
  OAI21_X1 U5110 ( .B1(n6110), .B2(n2945), .A(n4151), .ZN(U2857) );
  XNOR2_X1 U5111 ( .A(n4153), .B(n4152), .ZN(n6105) );
  AOI21_X1 U5112 ( .B1(n4156), .B2(n4155), .A(n4154), .ZN(n6160) );
  INV_X1 U5113 ( .A(n6160), .ZN(n4158) );
  INV_X1 U5114 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4157) );
  OAI22_X1 U5115 ( .A1(n5535), .A2(n4158), .B1(n4157), .B2(n5532), .ZN(n4159)
         );
  AOI21_X1 U5116 ( .B1(n6105), .B2(n5537), .A(n4159), .ZN(n4160) );
  INV_X1 U5117 ( .A(n4160), .ZN(U2856) );
  AOI22_X1 U5118 ( .A1(n6073), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6079), .ZN(n4162) );
  NAND2_X1 U5119 ( .A1(n4162), .A2(n4161), .ZN(U2940) );
  AOI22_X1 U5120 ( .A1(n6073), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n6079), .ZN(n4163) );
  INV_X1 U5121 ( .A(DATAI_13_), .ZN(n5126) );
  OR2_X1 U5122 ( .A1(n6058), .A2(n5126), .ZN(n4175) );
  NAND2_X1 U5123 ( .A1(n4163), .A2(n4175), .ZN(U2937) );
  AOI22_X1 U5124 ( .A1(n6073), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6079), .ZN(n4165) );
  NAND2_X1 U5125 ( .A1(n4165), .A2(n4164), .ZN(U2943) );
  AOI22_X1 U5126 ( .A1(n6073), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6079), .ZN(n4167) );
  NAND2_X1 U5127 ( .A1(n4167), .A2(n4166), .ZN(U2944) );
  AOI22_X1 U5128 ( .A1(n6073), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6079), .ZN(n4168) );
  NAND2_X1 U5129 ( .A1(n6080), .A2(DATAI_6_), .ZN(n4181) );
  NAND2_X1 U5130 ( .A1(n4168), .A2(n4181), .ZN(U2945) );
  AOI22_X1 U5131 ( .A1(n6073), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6079), .ZN(n4169) );
  NAND2_X1 U5132 ( .A1(n6080), .A2(DATAI_7_), .ZN(n4177) );
  NAND2_X1 U5133 ( .A1(n4169), .A2(n4177), .ZN(U2946) );
  AOI22_X1 U5134 ( .A1(n6073), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6079), .ZN(n4171) );
  NAND2_X1 U5135 ( .A1(n4171), .A2(n4170), .ZN(U2942) );
  AOI22_X1 U5136 ( .A1(n6073), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6079), .ZN(n4172) );
  NAND2_X1 U5137 ( .A1(n6080), .A2(DATAI_0_), .ZN(n4179) );
  NAND2_X1 U5138 ( .A1(n4172), .A2(n4179), .ZN(U2939) );
  AOI22_X1 U5139 ( .A1(n6073), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6079), .ZN(n4174) );
  NAND2_X1 U5140 ( .A1(n4174), .A2(n4173), .ZN(U2941) );
  AOI22_X1 U5141 ( .A1(n6073), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n6079), .ZN(n4176) );
  NAND2_X1 U5142 ( .A1(n4176), .A2(n4175), .ZN(U2952) );
  AOI22_X1 U5143 ( .A1(n6073), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6079), .ZN(n4178) );
  NAND2_X1 U5144 ( .A1(n4178), .A2(n4177), .ZN(U2931) );
  AOI22_X1 U5145 ( .A1(n6073), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6079), .ZN(n4180) );
  NAND2_X1 U5146 ( .A1(n4180), .A2(n4179), .ZN(U2924) );
  AOI22_X1 U5147 ( .A1(n6073), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6079), .ZN(n4182) );
  NAND2_X1 U5148 ( .A1(n4182), .A2(n4181), .ZN(U2930) );
  AOI22_X1 U5149 ( .A1(n6501), .A2(UWORD_REG_6__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4183) );
  OAI21_X1 U5150 ( .B1(n3765), .B2(n4195), .A(n4183), .ZN(U2901) );
  INV_X1 U5151 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4185) );
  AOI22_X1 U5152 ( .A1(n6501), .A2(UWORD_REG_4__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4184) );
  OAI21_X1 U5153 ( .B1(n4185), .B2(n4195), .A(n4184), .ZN(U2903) );
  INV_X1 U5154 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4187) );
  AOI22_X1 U5155 ( .A1(n6501), .A2(UWORD_REG_7__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4186) );
  OAI21_X1 U5156 ( .B1(n4187), .B2(n4195), .A(n4186), .ZN(U2900) );
  INV_X1 U5157 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4189) );
  AOI22_X1 U5158 ( .A1(n6501), .A2(UWORD_REG_5__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4188) );
  OAI21_X1 U5159 ( .B1(n4189), .B2(n4195), .A(n4188), .ZN(U2902) );
  AOI22_X1 U5160 ( .A1(n6501), .A2(UWORD_REG_3__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4190) );
  OAI21_X1 U5161 ( .B1(n3709), .B2(n4195), .A(n4190), .ZN(U2904) );
  AOI22_X1 U5162 ( .A1(n6041), .A2(UWORD_REG_1__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4191) );
  OAI21_X1 U5163 ( .B1(n3690), .B2(n4195), .A(n4191), .ZN(U2906) );
  INV_X1 U5164 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4193) );
  AOI22_X1 U5165 ( .A1(n6041), .A2(UWORD_REG_2__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4192) );
  OAI21_X1 U5166 ( .B1(n4193), .B2(n4195), .A(n4192), .ZN(U2905) );
  AOI22_X1 U5167 ( .A1(n6041), .A2(UWORD_REG_0__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4194) );
  OAI21_X1 U5168 ( .B1(n3652), .B2(n4195), .A(n4194), .ZN(U2907) );
  NAND2_X1 U5169 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5913), .ZN(n4222) );
  INV_X1 U5170 ( .A(n4222), .ZN(n4218) );
  NOR2_X1 U5171 ( .A1(n4196), .A2(n4232), .ZN(n4209) );
  NOR2_X1 U5172 ( .A1(n5152), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4197)
         );
  XNOR2_X1 U5173 ( .A(n4197), .B(n4206), .ZN(n4203) );
  XNOR2_X1 U5174 ( .A(n4198), .B(n4206), .ZN(n4201) );
  AOI21_X1 U5175 ( .B1(n5152), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n4206), 
        .ZN(n4199) );
  NOR2_X1 U5176 ( .A1(n3362), .A2(n4199), .ZN(n6485) );
  NOR2_X1 U5177 ( .A1(n4210), .A2(n6485), .ZN(n4200) );
  AOI21_X1 U5178 ( .B1(n6366), .B2(n4201), .A(n4200), .ZN(n4202) );
  OAI21_X1 U5179 ( .B1(n4209), .B2(n4203), .A(n4202), .ZN(n4204) );
  AOI21_X1 U5180 ( .B1(n6222), .B2(n4205), .A(n4204), .ZN(n6487) );
  MUX2_X1 U5181 ( .A(n6487), .B(n4206), .S(n6375), .Z(n6385) );
  INV_X1 U5182 ( .A(n5152), .ZN(n5392) );
  MUX2_X1 U5183 ( .A(n4210), .B(n4209), .S(n5392), .Z(n4208) );
  NAND2_X1 U5184 ( .A1(n6366), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4207) );
  NAND2_X1 U5185 ( .A1(n4208), .A2(n4207), .ZN(n4213) );
  MUX2_X1 U5186 ( .A(n4210), .B(n4209), .S(n5152), .Z(n4211) );
  NAND2_X1 U5187 ( .A1(n6366), .A2(n5404), .ZN(n5396) );
  NAND2_X1 U5188 ( .A1(n4211), .A2(n5396), .ZN(n4212) );
  MUX2_X1 U5189 ( .A(n4213), .B(n4212), .S(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .Z(n4214) );
  INV_X1 U5190 ( .A(n4214), .ZN(n4215) );
  OAI21_X1 U5191 ( .B1(n5397), .B2(n4894), .A(n4215), .ZN(n5155) );
  NAND2_X1 U5192 ( .A1(n6375), .A2(n5157), .ZN(n4216) );
  OAI21_X1 U5193 ( .B1(n5155), .B2(n6375), .A(n4216), .ZN(n6380) );
  NOR3_X1 U5194 ( .A1(n6385), .A2(STATE2_REG_1__SCAN_IN), .A3(n6380), .ZN(
        n4217) );
  AOI21_X1 U5195 ( .B1(n4219), .B2(n4218), .A(n4217), .ZN(n6386) );
  NOR2_X1 U5196 ( .A1(n6386), .A2(n5391), .ZN(n4229) );
  INV_X1 U5197 ( .A(n6309), .ZN(n4479) );
  NOR2_X1 U5198 ( .A1(n4220), .A2(n4479), .ZN(n4221) );
  XNOR2_X1 U5199 ( .A(n4221), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4609)
         );
  INV_X1 U5200 ( .A(n4609), .ZN(n5902) );
  INV_X1 U5201 ( .A(n4243), .ZN(n5901) );
  AOI22_X1 U5202 ( .A1(n5902), .A2(n5901), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6375), .ZN(n4223) );
  OAI22_X1 U5203 ( .A1(n4223), .A2(STATE2_REG_1__SCAN_IN), .B1(n4222), .B2(
        n6607), .ZN(n6392) );
  NOR3_X1 U5204 ( .A1(n4229), .A2(n6392), .A3(FLUSH_REG_SCAN_IN), .ZN(n4224)
         );
  OAI21_X1 U5205 ( .B1(n4224), .B2(n6480), .A(n5757), .ZN(n6182) );
  AND2_X1 U5206 ( .A1(n4554), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6186) );
  INV_X1 U5207 ( .A(n6186), .ZN(n6254) );
  NAND2_X1 U5208 ( .A1(n4614), .A2(n6186), .ZN(n5697) );
  NAND2_X1 U5209 ( .A1(n5697), .A2(n6500), .ZN(n5701) );
  AOI21_X1 U5210 ( .B1(n6187), .B2(n6254), .A(n5701), .ZN(n4226) );
  NAND2_X1 U5211 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6483), .ZN(n5699) );
  INV_X1 U5212 ( .A(n5699), .ZN(n5694) );
  NOR2_X1 U5213 ( .A1(n4894), .A2(n5694), .ZN(n4225) );
  OAI21_X1 U5214 ( .B1(n4226), .B2(n4225), .A(n6182), .ZN(n4227) );
  OAI21_X1 U5215 ( .B1(n6182), .B2(n6376), .A(n4227), .ZN(U3463) );
  NOR3_X1 U5216 ( .A1(n4229), .A2(n4228), .A3(n6392), .ZN(n6401) );
  OAI22_X1 U5217 ( .A1(n4615), .A2(n6308), .B1(n4654), .B2(n5694), .ZN(n4230)
         );
  OAI21_X1 U5218 ( .B1(n6401), .B2(n4230), .A(n6182), .ZN(n4231) );
  OAI21_X1 U5219 ( .B1(n6182), .B2(n4761), .A(n4231), .ZN(U3465) );
  INV_X1 U5220 ( .A(n6105), .ZN(n4250) );
  OR2_X1 U5221 ( .A1(n6407), .A2(n4234), .ZN(n4242) );
  INV_X1 U5222 ( .A(n4235), .ZN(n4241) );
  NAND4_X1 U5223 ( .A1(n4239), .A2(n4238), .A3(n4237), .A4(n4236), .ZN(n4240)
         );
  OAI22_X1 U5224 ( .A1(n4243), .A2(n4242), .B1(n4241), .B2(n4240), .ZN(n4244)
         );
  NOR2_X1 U5225 ( .A1(n4245), .A2(n4244), .ZN(n4246) );
  OR2_X1 U5226 ( .A1(n4247), .A2(n5422), .ZN(n4248) );
  AOI22_X1 U5227 ( .A1(n5544), .A2(DATAI_3_), .B1(EAX_REG_3__SCAN_IN), .B2(
        n6014), .ZN(n4249) );
  OAI21_X1 U5228 ( .B1(n4250), .B2(n5862), .A(n4249), .ZN(U2888) );
  OAI21_X1 U5229 ( .B1(n4251), .B2(n4256), .A(n4669), .ZN(n4472) );
  OAI21_X1 U5230 ( .B1(n4259), .B2(n4260), .A(n4252), .ZN(n4253) );
  NAND2_X1 U5231 ( .A1(n4253), .A2(n4595), .ZN(n4478) );
  OAI222_X1 U5232 ( .A1(n4472), .A2(n5535), .B1(n5532), .B2(n4469), .C1(n2945), 
        .C2(n4478), .ZN(U2853) );
  NAND2_X1 U5233 ( .A1(n4255), .A2(n4254), .ZN(n4258) );
  INV_X1 U5234 ( .A(n4256), .ZN(n4257) );
  NAND2_X1 U5235 ( .A1(n4258), .A2(n4257), .ZN(n6145) );
  XOR2_X1 U5236 ( .A(n4260), .B(n4259), .Z(n6097) );
  INV_X1 U5237 ( .A(n6097), .ZN(n4310) );
  OAI222_X1 U5238 ( .A1(n6145), .A2(n5535), .B1(n5532), .B2(n3007), .C1(n2945), 
        .C2(n4310), .ZN(U2854) );
  INV_X1 U5239 ( .A(DATAI_2_), .ZN(n6597) );
  INV_X1 U5240 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6037) );
  OAI222_X1 U5241 ( .A1(n6110), .A2(n5862), .B1(n5127), .B2(n6597), .C1(n5421), 
        .C2(n6037), .ZN(U2889) );
  INV_X1 U5242 ( .A(DATAI_4_), .ZN(n4264) );
  INV_X1 U5243 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6034) );
  OAI222_X1 U5244 ( .A1(n4664), .A2(n5862), .B1(n5127), .B2(n4264), .C1(n5421), 
        .C2(n6034), .ZN(U2887) );
  NOR2_X1 U5245 ( .A1(n4300), .A2(n4262), .ZN(n6338) );
  INV_X1 U5246 ( .A(n6338), .ZN(n4876) );
  NAND2_X1 U5247 ( .A1(n2946), .A2(DATAI_28_), .ZN(n6342) );
  INV_X1 U5248 ( .A(n6342), .ZN(n6278) );
  NAND2_X1 U5249 ( .A1(n4554), .A2(n4615), .ZN(n4831) );
  INV_X1 U5250 ( .A(n4831), .ZN(n4263) );
  AND2_X1 U5251 ( .A1(n4614), .A2(n4263), .ZN(n4485) );
  AND2_X1 U5252 ( .A1(n4485), .A2(n5696), .ZN(n4416) );
  INV_X1 U5253 ( .A(n6184), .ZN(n6252) );
  NOR3_X1 U5254 ( .A1(n6187), .A2(n4486), .A3(n6252), .ZN(n5703) );
  NAND2_X1 U5255 ( .A1(n2946), .A2(DATAI_20_), .ZN(n6281) );
  NAND2_X1 U5256 ( .A1(n6222), .A2(n6256), .ZN(n4311) );
  INV_X1 U5257 ( .A(n4886), .ZN(n5693) );
  OR2_X1 U5258 ( .A1(n4894), .A2(n5693), .ZN(n4621) );
  OAI21_X1 U5259 ( .B1(n4311), .B2(n4621), .A(n4306), .ZN(n4268) );
  AOI22_X1 U5260 ( .A1(n4268), .A2(n6500), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4272), .ZN(n4301) );
  NOR2_X1 U5261 ( .A1(n4264), .A2(n5757), .ZN(n6337) );
  INV_X1 U5262 ( .A(n6337), .ZN(n5783) );
  OAI22_X1 U5263 ( .A1(n5743), .A2(n6281), .B1(n4301), .B2(n5783), .ZN(n4265)
         );
  AOI21_X1 U5264 ( .B1(n6278), .B2(n4416), .A(n4265), .ZN(n4274) );
  INV_X1 U5265 ( .A(n4554), .ZN(n4525) );
  NOR3_X1 U5266 ( .A1(n6187), .A2(n4486), .A3(n4525), .ZN(n4267) );
  NOR2_X1 U5267 ( .A1(n6308), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6224) );
  INV_X1 U5268 ( .A(n6224), .ZN(n5752) );
  OAI21_X1 U5269 ( .B1(n4267), .B2(n5591), .A(n5752), .ZN(n4270) );
  INV_X1 U5270 ( .A(n4268), .ZN(n4269) );
  NAND2_X1 U5271 ( .A1(n4270), .A2(n4269), .ZN(n4271) );
  OAI211_X1 U5272 ( .C1(n6500), .C2(n4272), .A(n4271), .B(n6259), .ZN(n4303)
         );
  NAND2_X1 U5273 ( .A1(n4303), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4273)
         );
  OAI211_X1 U5274 ( .C1(n4876), .C2(n4306), .A(n4274), .B(n4273), .ZN(U3144)
         );
  NOR2_X1 U5275 ( .A1(n4300), .A2(n4275), .ZN(n6344) );
  INV_X1 U5276 ( .A(n6344), .ZN(n4852) );
  NAND2_X1 U5277 ( .A1(n2946), .A2(DATAI_29_), .ZN(n6348) );
  INV_X1 U5278 ( .A(n6348), .ZN(n6282) );
  NAND2_X1 U5279 ( .A1(n2946), .A2(DATAI_21_), .ZN(n6285) );
  NOR2_X1 U5280 ( .A1(n4276), .A2(n5757), .ZN(n6343) );
  INV_X1 U5281 ( .A(n6343), .ZN(n5788) );
  OAI22_X1 U5282 ( .A1(n5743), .A2(n6285), .B1(n4301), .B2(n5788), .ZN(n4277)
         );
  AOI21_X1 U5283 ( .B1(n6282), .B2(n4416), .A(n4277), .ZN(n4279) );
  NAND2_X1 U5284 ( .A1(n4303), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4278)
         );
  OAI211_X1 U5285 ( .C1(n4852), .C2(n4306), .A(n4279), .B(n4278), .ZN(U3145)
         );
  NOR2_X1 U5286 ( .A1(n4300), .A2(n4280), .ZN(n6326) );
  INV_X1 U5287 ( .A(n6326), .ZN(n4848) );
  NAND2_X1 U5288 ( .A1(n2946), .A2(DATAI_26_), .ZN(n6330) );
  INV_X1 U5289 ( .A(n6330), .ZN(n6270) );
  NAND2_X1 U5290 ( .A1(n2946), .A2(DATAI_18_), .ZN(n6273) );
  NOR2_X1 U5291 ( .A1(n6597), .A2(n5757), .ZN(n6325) );
  INV_X1 U5292 ( .A(n6325), .ZN(n5773) );
  OAI22_X1 U5293 ( .A1(n5743), .A2(n6273), .B1(n4301), .B2(n5773), .ZN(n4281)
         );
  AOI21_X1 U5294 ( .B1(n6270), .B2(n4416), .A(n4281), .ZN(n4283) );
  NAND2_X1 U5295 ( .A1(n4303), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4282)
         );
  OAI211_X1 U5296 ( .C1(n4848), .C2(n4306), .A(n4283), .B(n4282), .ZN(U3142)
         );
  NOR2_X1 U5297 ( .A1(n4300), .A2(n4284), .ZN(n6320) );
  INV_X1 U5298 ( .A(n6320), .ZN(n4860) );
  NAND2_X1 U5299 ( .A1(n2946), .A2(DATAI_25_), .ZN(n6324) );
  INV_X1 U5300 ( .A(n6324), .ZN(n6266) );
  NAND2_X1 U5301 ( .A1(n2946), .A2(DATAI_17_), .ZN(n6269) );
  INV_X1 U5302 ( .A(DATAI_1_), .ZN(n4307) );
  NOR2_X1 U5303 ( .A1(n4307), .A2(n5757), .ZN(n6319) );
  INV_X1 U5304 ( .A(n6319), .ZN(n5768) );
  OAI22_X1 U5305 ( .A1(n5743), .A2(n6269), .B1(n4301), .B2(n5768), .ZN(n4285)
         );
  AOI21_X1 U5306 ( .B1(n6266), .B2(n4416), .A(n4285), .ZN(n4287) );
  NAND2_X1 U5307 ( .A1(n4303), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4286)
         );
  OAI211_X1 U5308 ( .C1(n4860), .C2(n4306), .A(n4287), .B(n4286), .ZN(U3141)
         );
  NOR2_X1 U5309 ( .A1(n4300), .A2(n4288), .ZN(n6332) );
  INV_X1 U5310 ( .A(n6332), .ZN(n4844) );
  NAND2_X1 U5311 ( .A1(n2946), .A2(DATAI_27_), .ZN(n6336) );
  INV_X1 U5312 ( .A(n6336), .ZN(n6274) );
  NAND2_X1 U5313 ( .A1(n2946), .A2(DATAI_19_), .ZN(n6277) );
  INV_X1 U5314 ( .A(DATAI_3_), .ZN(n6625) );
  NOR2_X1 U5315 ( .A1(n6625), .A2(n5757), .ZN(n6331) );
  INV_X1 U5316 ( .A(n6331), .ZN(n5778) );
  OAI22_X1 U5317 ( .A1(n5743), .A2(n6277), .B1(n4301), .B2(n5778), .ZN(n4289)
         );
  AOI21_X1 U5318 ( .B1(n6274), .B2(n4416), .A(n4289), .ZN(n4291) );
  NAND2_X1 U5319 ( .A1(n4303), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4290)
         );
  OAI211_X1 U5320 ( .C1(n4844), .C2(n4306), .A(n4291), .B(n4290), .ZN(U3143)
         );
  NOR2_X1 U5321 ( .A1(n4300), .A2(n4292), .ZN(n6350) );
  INV_X1 U5322 ( .A(n6350), .ZN(n4856) );
  NAND2_X1 U5323 ( .A1(n2946), .A2(DATAI_30_), .ZN(n6354) );
  INV_X1 U5324 ( .A(n6354), .ZN(n6286) );
  NAND2_X1 U5325 ( .A1(n2946), .A2(DATAI_22_), .ZN(n6290) );
  INV_X1 U5326 ( .A(DATAI_6_), .ZN(n4308) );
  NOR2_X1 U5327 ( .A1(n4308), .A2(n5757), .ZN(n6349) );
  INV_X1 U5328 ( .A(n6349), .ZN(n5793) );
  OAI22_X1 U5329 ( .A1(n5743), .A2(n6290), .B1(n4301), .B2(n5793), .ZN(n4293)
         );
  AOI21_X1 U5330 ( .B1(n6286), .B2(n4416), .A(n4293), .ZN(n4295) );
  NAND2_X1 U5331 ( .A1(n4303), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4294)
         );
  OAI211_X1 U5332 ( .C1(n4856), .C2(n4306), .A(n4295), .B(n4294), .ZN(U3146)
         );
  NOR2_X1 U5333 ( .A1(n4300), .A2(n5422), .ZN(n6358) );
  INV_X1 U5334 ( .A(n6358), .ZN(n4868) );
  NAND2_X1 U5335 ( .A1(n2946), .A2(DATAI_31_), .ZN(n6365) );
  INV_X1 U5336 ( .A(n6365), .ZN(n6211) );
  NAND2_X1 U5337 ( .A1(n2946), .A2(DATAI_23_), .ZN(n6218) );
  INV_X1 U5338 ( .A(DATAI_7_), .ZN(n4597) );
  NOR2_X1 U5339 ( .A1(n4597), .A2(n5757), .ZN(n6356) );
  INV_X1 U5340 ( .A(n6356), .ZN(n5798) );
  OAI22_X1 U5341 ( .A1(n5743), .A2(n6218), .B1(n4301), .B2(n5798), .ZN(n4296)
         );
  AOI21_X1 U5342 ( .B1(n6211), .B2(n4416), .A(n4296), .ZN(n4298) );
  NAND2_X1 U5343 ( .A1(n4303), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4297)
         );
  OAI211_X1 U5344 ( .C1(n4868), .C2(n4306), .A(n4298), .B(n4297), .ZN(U3147)
         );
  NOR2_X1 U5345 ( .A1(n4300), .A2(n4299), .ZN(n6304) );
  INV_X1 U5346 ( .A(n6304), .ZN(n4864) );
  NAND2_X1 U5347 ( .A1(n2946), .A2(DATAI_24_), .ZN(n6318) );
  INV_X1 U5348 ( .A(n6318), .ZN(n6185) );
  NAND2_X1 U5349 ( .A1(n2946), .A2(DATAI_16_), .ZN(n6198) );
  INV_X1 U5350 ( .A(DATAI_0_), .ZN(n6549) );
  NOR2_X1 U5351 ( .A1(n6549), .A2(n5757), .ZN(n6303) );
  INV_X1 U5352 ( .A(n6303), .ZN(n5762) );
  OAI22_X1 U5353 ( .A1(n5743), .A2(n6198), .B1(n4301), .B2(n5762), .ZN(n4302)
         );
  AOI21_X1 U5354 ( .B1(n6185), .B2(n4416), .A(n4302), .ZN(n4305) );
  NAND2_X1 U5355 ( .A1(n4303), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4304)
         );
  OAI211_X1 U5356 ( .C1(n4864), .C2(n4306), .A(n4305), .B(n4304), .ZN(U3140)
         );
  INV_X1 U5357 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6039) );
  OAI222_X1 U5358 ( .A1(n4889), .A2(n5862), .B1(n5127), .B2(n4307), .C1(n5421), 
        .C2(n6039), .ZN(U2890) );
  INV_X1 U5359 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6537) );
  OAI222_X1 U5360 ( .A1(n4478), .A2(n5862), .B1(n5127), .B2(n4308), .C1(n5421), 
        .C2(n6537), .ZN(U2885) );
  INV_X1 U5361 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6044) );
  OAI222_X1 U5362 ( .A1(n4659), .A2(n5862), .B1(n5127), .B2(n6549), .C1(n5421), 
        .C2(n6044), .ZN(U2891) );
  OAI222_X1 U5363 ( .A1(n5127), .A2(n4276), .B1(n5862), .B2(n4310), .C1(n4309), 
        .C2(n5421), .ZN(U2886) );
  NOR2_X1 U5364 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6376), .ZN(n4760)
         );
  NAND2_X1 U5365 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4760), .ZN(n6298) );
  NOR2_X1 U5366 ( .A1(n4761), .A2(n6298), .ZN(n4312) );
  INV_X1 U5367 ( .A(n4312), .ZN(n4341) );
  INV_X1 U5368 ( .A(n4311), .ZN(n4553) );
  OR2_X1 U5369 ( .A1(n4894), .A2(n4886), .ZN(n6223) );
  INV_X1 U5370 ( .A(n6223), .ZN(n6310) );
  AOI21_X1 U5371 ( .B1(n4553), .B2(n6310), .A(n4312), .ZN(n4320) );
  NOR2_X1 U5372 ( .A1(n4486), .A2(n4554), .ZN(n4313) );
  NAND2_X1 U5373 ( .A1(n4614), .A2(n4313), .ZN(n4321) );
  OR2_X1 U5374 ( .A1(n4321), .A2(n6305), .ZN(n4314) );
  AND2_X1 U5375 ( .A1(n4314), .A2(n6500), .ZN(n4316) );
  AOI22_X1 U5376 ( .A1(n4320), .A2(n4316), .B1(n6308), .B2(n6298), .ZN(n4315)
         );
  NAND2_X1 U5377 ( .A1(n6259), .A2(n4315), .ZN(n4338) );
  INV_X1 U5378 ( .A(n4316), .ZN(n4319) );
  INV_X1 U5379 ( .A(n4760), .ZN(n4318) );
  NAND2_X1 U5380 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4317) );
  OAI22_X1 U5381 ( .A1(n4320), .A2(n4319), .B1(n4318), .B2(n4317), .ZN(n4337)
         );
  AOI22_X1 U5382 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4338), .B1(n6303), 
        .B2(n4337), .ZN(n4324) );
  INV_X1 U5383 ( .A(n6198), .ZN(n6315) );
  NOR2_X2 U5384 ( .A1(n4321), .A2(n4615), .ZN(n4445) );
  INV_X1 U5385 ( .A(n4321), .ZN(n4322) );
  AOI22_X1 U5386 ( .A1(n6315), .A2(n4445), .B1(n6359), .B2(n6185), .ZN(n4323)
         );
  OAI211_X1 U5387 ( .C1(n4864), .C2(n4341), .A(n4324), .B(n4323), .ZN(U3124)
         );
  AOI22_X1 U5388 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4338), .B1(n6337), 
        .B2(n4337), .ZN(n4326) );
  INV_X1 U5389 ( .A(n6281), .ZN(n6339) );
  AOI22_X1 U5390 ( .A1(n6339), .A2(n4445), .B1(n6359), .B2(n6278), .ZN(n4325)
         );
  OAI211_X1 U5391 ( .C1(n4876), .C2(n4341), .A(n4326), .B(n4325), .ZN(U3128)
         );
  AOI22_X1 U5392 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4338), .B1(n6319), 
        .B2(n4337), .ZN(n4328) );
  INV_X1 U5393 ( .A(n6269), .ZN(n6321) );
  AOI22_X1 U5394 ( .A1(n6321), .A2(n4445), .B1(n6359), .B2(n6266), .ZN(n4327)
         );
  OAI211_X1 U5395 ( .C1(n4860), .C2(n4341), .A(n4328), .B(n4327), .ZN(U3125)
         );
  AOI22_X1 U5396 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4338), .B1(n6349), 
        .B2(n4337), .ZN(n4330) );
  INV_X1 U5397 ( .A(n6290), .ZN(n6351) );
  AOI22_X1 U5398 ( .A1(n6351), .A2(n4445), .B1(n6359), .B2(n6286), .ZN(n4329)
         );
  OAI211_X1 U5399 ( .C1(n4856), .C2(n4341), .A(n4330), .B(n4329), .ZN(U3130)
         );
  AOI22_X1 U5400 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4338), .B1(n6343), 
        .B2(n4337), .ZN(n4332) );
  INV_X1 U5401 ( .A(n6285), .ZN(n6345) );
  AOI22_X1 U5402 ( .A1(n6345), .A2(n4445), .B1(n6359), .B2(n6282), .ZN(n4331)
         );
  OAI211_X1 U5403 ( .C1(n4852), .C2(n4341), .A(n4332), .B(n4331), .ZN(U3129)
         );
  AOI22_X1 U5404 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4338), .B1(n6331), 
        .B2(n4337), .ZN(n4334) );
  INV_X1 U5405 ( .A(n6277), .ZN(n6333) );
  AOI22_X1 U5406 ( .A1(n6333), .A2(n4445), .B1(n6359), .B2(n6274), .ZN(n4333)
         );
  OAI211_X1 U5407 ( .C1(n4844), .C2(n4341), .A(n4334), .B(n4333), .ZN(U3127)
         );
  AOI22_X1 U5408 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4338), .B1(n6325), 
        .B2(n4337), .ZN(n4336) );
  INV_X1 U5409 ( .A(n6273), .ZN(n6327) );
  AOI22_X1 U5410 ( .A1(n6327), .A2(n4445), .B1(n6359), .B2(n6270), .ZN(n4335)
         );
  OAI211_X1 U5411 ( .C1(n4848), .C2(n4341), .A(n4336), .B(n4335), .ZN(U3126)
         );
  AOI22_X1 U5412 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4338), .B1(n6356), 
        .B2(n4337), .ZN(n4340) );
  INV_X1 U5413 ( .A(n6218), .ZN(n6360) );
  AOI22_X1 U5414 ( .A1(n6360), .A2(n4445), .B1(n6359), .B2(n6211), .ZN(n4339)
         );
  OAI211_X1 U5415 ( .C1(n4868), .C2(n4341), .A(n4340), .B(n4339), .ZN(U3131)
         );
  NAND2_X1 U5416 ( .A1(n4832), .A2(n4676), .ZN(n4345) );
  NAND2_X1 U5417 ( .A1(n4354), .A2(n4353), .ZN(n4352) );
  NAND2_X1 U5418 ( .A1(n4352), .A2(n4347), .ZN(n4373) );
  INV_X1 U5419 ( .A(n4372), .ZN(n4342) );
  XNOR2_X1 U5420 ( .A(n4373), .B(n4342), .ZN(n4343) );
  NAND2_X1 U5421 ( .A1(n4343), .A2(n4697), .ZN(n4344) );
  NAND2_X1 U5422 ( .A1(n4345), .A2(n4344), .ZN(n4369) );
  INV_X1 U5423 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6165) );
  XNOR2_X1 U5424 ( .A(n4369), .B(n6165), .ZN(n6102) );
  NAND2_X1 U5425 ( .A1(n4346), .A2(n4676), .ZN(n4351) );
  XNOR2_X1 U5426 ( .A(n4352), .B(n4347), .ZN(n4349) );
  AOI21_X1 U5427 ( .B1(n4349), .B2(n4697), .A(n4348), .ZN(n4350) );
  NAND2_X1 U5428 ( .A1(n4351), .A2(n4350), .ZN(n6112) );
  NAND2_X1 U5429 ( .A1(n6112), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4366)
         );
  NAND2_X1 U5430 ( .A1(n4266), .A2(n4676), .ZN(n4359) );
  OAI21_X1 U5431 ( .B1(n4354), .B2(n4353), .A(n4352), .ZN(n4356) );
  OAI211_X1 U5432 ( .C1(n4356), .C2(n6506), .A(n3263), .B(n5190), .ZN(n4357)
         );
  INV_X1 U5433 ( .A(n4357), .ZN(n4358) );
  NAND2_X1 U5434 ( .A1(n4359), .A2(n4358), .ZN(n4406) );
  NAND2_X1 U5435 ( .A1(n4362), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4360)
         );
  INV_X1 U5436 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6583) );
  NAND2_X1 U5437 ( .A1(n4360), .A2(n6583), .ZN(n4363) );
  AND2_X1 U5438 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4361) );
  NAND2_X1 U5439 ( .A1(n4362), .A2(n4361), .ZN(n4364) );
  AND2_X1 U5440 ( .A1(n4363), .A2(n4364), .ZN(n4405) );
  INV_X1 U5441 ( .A(n4364), .ZN(n4365) );
  NAND2_X1 U5442 ( .A1(n4366), .A2(n6111), .ZN(n4368) );
  OR2_X1 U5443 ( .A1(n6112), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4367)
         );
  AND2_X1 U5444 ( .A1(n4368), .A2(n4367), .ZN(n6101) );
  NAND2_X1 U5445 ( .A1(n6102), .A2(n6101), .ZN(n6103) );
  NAND2_X1 U5446 ( .A1(n4369), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4370)
         );
  NAND2_X1 U5447 ( .A1(n6103), .A2(n4370), .ZN(n4662) );
  NAND2_X1 U5448 ( .A1(n4371), .A2(n4676), .ZN(n4376) );
  NAND2_X1 U5449 ( .A1(n4373), .A2(n4372), .ZN(n4392) );
  XNOR2_X1 U5450 ( .A(n4392), .B(n4389), .ZN(n4374) );
  NAND2_X1 U5451 ( .A1(n4374), .A2(n4697), .ZN(n4375) );
  NAND2_X1 U5452 ( .A1(n4376), .A2(n4375), .ZN(n4377) );
  XNOR2_X1 U5453 ( .A(n4377), .B(n6159), .ZN(n4661) );
  NAND2_X1 U5454 ( .A1(n4662), .A2(n4661), .ZN(n4660) );
  NAND2_X1 U5455 ( .A1(n4377), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4378)
         );
  NAND2_X1 U5456 ( .A1(n4660), .A2(n4378), .ZN(n6095) );
  NAND2_X1 U5457 ( .A1(n4379), .A2(n4676), .ZN(n4384) );
  INV_X1 U5458 ( .A(n4389), .ZN(n4380) );
  OR2_X1 U5459 ( .A1(n4392), .A2(n4380), .ZN(n4381) );
  XNOR2_X1 U5460 ( .A(n4381), .B(n4390), .ZN(n4382) );
  NAND2_X1 U5461 ( .A1(n4382), .A2(n4697), .ZN(n4383) );
  NAND2_X1 U5462 ( .A1(n4384), .A2(n4383), .ZN(n4386) );
  INV_X1 U5463 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4385) );
  XNOR2_X1 U5464 ( .A(n4386), .B(n4385), .ZN(n6094) );
  NAND2_X1 U5465 ( .A1(n6095), .A2(n6094), .ZN(n6093) );
  NAND2_X1 U5466 ( .A1(n4386), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4387)
         );
  NAND2_X1 U5467 ( .A1(n6093), .A2(n4387), .ZN(n4688) );
  NAND3_X1 U5468 ( .A1(n4694), .A2(n4388), .A3(n4676), .ZN(n4395) );
  NAND2_X1 U5469 ( .A1(n4390), .A2(n4389), .ZN(n4391) );
  OR2_X1 U5470 ( .A1(n4392), .A2(n4391), .ZN(n4678) );
  XNOR2_X1 U5471 ( .A(n4678), .B(n4679), .ZN(n4393) );
  NAND2_X1 U5472 ( .A1(n4393), .A2(n4697), .ZN(n4394) );
  NAND2_X1 U5473 ( .A1(n4395), .A2(n4394), .ZN(n4685) );
  INV_X1 U5474 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4396) );
  XNOR2_X1 U5475 ( .A(n4685), .B(n4396), .ZN(n4684) );
  NAND2_X1 U5476 ( .A1(n4688), .A2(n4684), .ZN(n6084) );
  OAI21_X1 U5477 ( .B1(n4688), .B2(n4684), .A(n6084), .ZN(n4455) );
  INV_X1 U5478 ( .A(n4472), .ZN(n4403) );
  INV_X1 U5479 ( .A(REIP_REG_6__SCAN_IN), .ZN(n4397) );
  NOR2_X1 U5480 ( .A1(n5585), .A2(n4397), .ZN(n4449) );
  NOR2_X1 U5481 ( .A1(n6173), .A2(n6583), .ZN(n6176) );
  OR2_X1 U5482 ( .A1(n4965), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5686)
         );
  INV_X1 U5483 ( .A(n5074), .ZN(n6175) );
  AOI21_X1 U5484 ( .B1(n6176), .B2(n6174), .A(n6175), .ZN(n6155) );
  AOI21_X1 U5485 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6177) );
  NAND2_X1 U5486 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6156) );
  NOR2_X1 U5487 ( .A1(n6177), .A2(n6156), .ZN(n6144) );
  NAND2_X1 U5488 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6144), .ZN(n4399)
         );
  NOR2_X1 U5489 ( .A1(n6155), .A2(n4399), .ZN(n4401) );
  INV_X1 U5490 ( .A(n4965), .ZN(n4398) );
  NAND2_X1 U5491 ( .A1(n4967), .A2(n4398), .ZN(n5687) );
  INV_X1 U5492 ( .A(n5052), .ZN(n4818) );
  NAND2_X1 U5493 ( .A1(n5685), .A2(n5074), .ZN(n5054) );
  OAI21_X1 U5494 ( .B1(n4818), .B2(n6176), .A(n5054), .ZN(n6172) );
  AOI21_X1 U5495 ( .B1(n5687), .B2(n4399), .A(n6172), .ZN(n6151) );
  INV_X1 U5496 ( .A(n6151), .ZN(n4400) );
  MUX2_X1 U5497 ( .A(n4401), .B(n4400), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4402) );
  AOI211_X1 U5498 ( .C1(n6168), .C2(n4403), .A(n4449), .B(n4402), .ZN(n4404)
         );
  OAI21_X1 U5499 ( .B1(n5680), .B2(n4455), .A(n4404), .ZN(U3012) );
  XNOR2_X1 U5500 ( .A(n4406), .B(n4405), .ZN(n5681) );
  INV_X1 U5501 ( .A(n4889), .ZN(n4410) );
  INV_X1 U5502 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6490) );
  NOR2_X1 U5503 ( .A1(n5585), .A2(n6490), .ZN(n5683) );
  AOI21_X1 U5504 ( .B1(n6109), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n5683), 
        .ZN(n4408) );
  OAI21_X1 U5505 ( .B1(n6118), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4408), 
        .ZN(n4409) );
  AOI21_X1 U5506 ( .B1(n4410), .B2(n2946), .A(n4409), .ZN(n4411) );
  OAI21_X1 U5507 ( .B1(n5681), .B2(n5912), .A(n4411), .ZN(U2985) );
  OR2_X1 U5508 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4412), .ZN(n4448)
         );
  NOR3_X1 U5509 ( .A1(n4445), .A2(n4416), .A3(n6308), .ZN(n4413) );
  NOR2_X1 U5510 ( .A1(n4413), .A2(n6224), .ZN(n4415) );
  INV_X1 U5511 ( .A(n6222), .ZN(n6301) );
  NOR2_X1 U5512 ( .A1(n6301), .A2(n4621), .ZN(n4419) );
  NOR2_X1 U5513 ( .A1(n4417), .A2(n6405), .ZN(n6226) );
  OAI21_X1 U5514 ( .B1(n5756), .B2(n6405), .A(n5708), .ZN(n4727) );
  NOR2_X1 U5515 ( .A1(n6226), .A2(n4727), .ZN(n4618) );
  NOR2_X1 U5516 ( .A1(n6405), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4728)
         );
  AOI21_X1 U5517 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n4448), .A(n4728), .ZN(
        n4414) );
  OAI211_X1 U5518 ( .C1(n4415), .C2(n4419), .A(n4618), .B(n4414), .ZN(n4441)
         );
  NAND2_X1 U5519 ( .A1(n4441), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4422)
         );
  INV_X1 U5520 ( .A(n4416), .ZN(n4443) );
  AND2_X1 U5521 ( .A1(n4417), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5709) );
  INV_X1 U5522 ( .A(n5709), .ZN(n6300) );
  NOR2_X1 U5523 ( .A1(n6300), .A2(n6383), .ZN(n4418) );
  AOI22_X1 U5524 ( .A1(n4419), .A2(n6500), .B1(n5756), .B2(n4418), .ZN(n4442)
         );
  OAI22_X1 U5525 ( .A1(n4443), .A2(n6273), .B1(n4442), .B2(n5773), .ZN(n4420)
         );
  AOI21_X1 U5526 ( .B1(n6270), .B2(n4445), .A(n4420), .ZN(n4421) );
  OAI211_X1 U5527 ( .C1(n4448), .C2(n4848), .A(n4422), .B(n4421), .ZN(U3134)
         );
  NAND2_X1 U5528 ( .A1(n4441), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4425)
         );
  OAI22_X1 U5529 ( .A1(n4443), .A2(n6218), .B1(n4442), .B2(n5798), .ZN(n4423)
         );
  AOI21_X1 U5530 ( .B1(n6211), .B2(n4445), .A(n4423), .ZN(n4424) );
  OAI211_X1 U5531 ( .C1(n4448), .C2(n4868), .A(n4425), .B(n4424), .ZN(U3139)
         );
  NAND2_X1 U5532 ( .A1(n4441), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4428)
         );
  OAI22_X1 U5533 ( .A1(n4443), .A2(n6281), .B1(n4442), .B2(n5783), .ZN(n4426)
         );
  AOI21_X1 U5534 ( .B1(n6278), .B2(n4445), .A(n4426), .ZN(n4427) );
  OAI211_X1 U5535 ( .C1(n4448), .C2(n4876), .A(n4428), .B(n4427), .ZN(U3136)
         );
  NAND2_X1 U5536 ( .A1(n4441), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4431)
         );
  OAI22_X1 U5537 ( .A1(n4443), .A2(n6269), .B1(n4442), .B2(n5768), .ZN(n4429)
         );
  AOI21_X1 U5538 ( .B1(n6266), .B2(n4445), .A(n4429), .ZN(n4430) );
  OAI211_X1 U5539 ( .C1(n4448), .C2(n4860), .A(n4431), .B(n4430), .ZN(U3133)
         );
  NAND2_X1 U5540 ( .A1(n4441), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4434)
         );
  OAI22_X1 U5541 ( .A1(n4443), .A2(n6285), .B1(n4442), .B2(n5788), .ZN(n4432)
         );
  AOI21_X1 U5542 ( .B1(n6282), .B2(n4445), .A(n4432), .ZN(n4433) );
  OAI211_X1 U5543 ( .C1(n4448), .C2(n4852), .A(n4434), .B(n4433), .ZN(U3137)
         );
  NAND2_X1 U5544 ( .A1(n4441), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4437)
         );
  OAI22_X1 U5545 ( .A1(n4443), .A2(n6277), .B1(n4442), .B2(n5778), .ZN(n4435)
         );
  AOI21_X1 U5546 ( .B1(n6274), .B2(n4445), .A(n4435), .ZN(n4436) );
  OAI211_X1 U5547 ( .C1(n4448), .C2(n4844), .A(n4437), .B(n4436), .ZN(U3135)
         );
  NAND2_X1 U5548 ( .A1(n4441), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4440)
         );
  OAI22_X1 U5549 ( .A1(n4443), .A2(n6198), .B1(n4442), .B2(n5762), .ZN(n4438)
         );
  AOI21_X1 U5550 ( .B1(n6185), .B2(n4445), .A(n4438), .ZN(n4439) );
  OAI211_X1 U5551 ( .C1(n4864), .C2(n4448), .A(n4440), .B(n4439), .ZN(U3132)
         );
  NAND2_X1 U5552 ( .A1(n4441), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4447)
         );
  OAI22_X1 U5553 ( .A1(n4443), .A2(n6290), .B1(n4442), .B2(n5793), .ZN(n4444)
         );
  AOI21_X1 U5554 ( .B1(n6286), .B2(n4445), .A(n4444), .ZN(n4446) );
  OAI211_X1 U5555 ( .C1(n4448), .C2(n4856), .A(n4447), .B(n4446), .ZN(U3138)
         );
  INV_X1 U5556 ( .A(n4478), .ZN(n4453) );
  INV_X1 U5557 ( .A(n4475), .ZN(n4451) );
  AOI21_X1 U5558 ( .B1(n6109), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n4449), 
        .ZN(n4450) );
  OAI21_X1 U5559 ( .B1(n6118), .B2(n4451), .A(n4450), .ZN(n4452) );
  AOI21_X1 U5560 ( .B1(n4453), .B2(n2946), .A(n4452), .ZN(n4454) );
  OAI21_X1 U5561 ( .B1(n4455), .B2(n5912), .A(n4454), .ZN(U2980) );
  INV_X1 U5562 ( .A(n4456), .ZN(n4457) );
  NAND2_X1 U5563 ( .A1(n4992), .A2(n4457), .ZN(n4458) );
  NAND2_X1 U5564 ( .A1(n5459), .A2(n4458), .ZN(n5986) );
  INV_X1 U5565 ( .A(n5979), .ZN(n4460) );
  INV_X1 U5566 ( .A(REIP_REG_5__SCAN_IN), .ZN(n4459) );
  OR3_X1 U5567 ( .A1(n5978), .A2(n4460), .A3(n4459), .ZN(n5973) );
  AOI22_X1 U5568 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5986), .B1(n5973), .B2(n4397), .ZN(n4461) );
  INV_X1 U5569 ( .A(n4461), .ZN(n4477) );
  INV_X1 U5570 ( .A(n4462), .ZN(n4463) );
  NAND2_X1 U5571 ( .A1(n4697), .A2(n6399), .ZN(n4467) );
  INV_X1 U5572 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5412) );
  NAND3_X1 U5573 ( .A1(n3187), .A2(n5412), .A3(n4464), .ZN(n4466) );
  NAND2_X1 U5574 ( .A1(n4467), .A2(n4466), .ZN(n4468) );
  AND2_X2 U5575 ( .A1(n4602), .A2(n4468), .ZN(n5993) );
  INV_X1 U5576 ( .A(n5993), .ZN(n5954) );
  NOR2_X1 U5577 ( .A1(n5954), .A2(n4469), .ZN(n4474) );
  NAND2_X1 U5578 ( .A1(n4992), .A2(n4470), .ZN(n5982) );
  NAND2_X1 U5579 ( .A1(n5991), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4471)
         );
  OAI211_X1 U5580 ( .C1(n5983), .C2(n4472), .A(n5982), .B(n4471), .ZN(n4473)
         );
  AOI211_X1 U5581 ( .C1(n5958), .C2(n4475), .A(n4474), .B(n4473), .ZN(n4476)
         );
  OAI211_X1 U5582 ( .C1(n4478), .C2(n5820), .A(n4477), .B(n4476), .ZN(U2821)
         );
  OAI21_X1 U5583 ( .B1(n4486), .B2(n6308), .A(n5701), .ZN(n4483) );
  NAND2_X1 U5584 ( .A1(n6256), .A2(n4479), .ZN(n4763) );
  OAI21_X1 U5585 ( .B1(n4621), .B2(n4763), .A(n4517), .ZN(n4482) );
  INV_X1 U5586 ( .A(n4482), .ZN(n4481) );
  OAI21_X1 U5587 ( .B1(n6500), .B2(n4612), .A(n6259), .ZN(n4480) );
  AOI21_X1 U5588 ( .B1(n4483), .B2(n4481), .A(n4480), .ZN(n4522) );
  INV_X1 U5589 ( .A(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4491) );
  AOI22_X1 U5590 ( .A1(n4483), .A2(n4482), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4612), .ZN(n4484) );
  AND2_X1 U5591 ( .A1(n6184), .A2(n4486), .ZN(n4487) );
  NAND2_X1 U5592 ( .A1(n4614), .A2(n4487), .ZN(n5800) );
  INV_X1 U5593 ( .A(n5800), .ZN(n4515) );
  AOI22_X1 U5594 ( .A1(n4620), .A2(n6274), .B1(n6333), .B2(n4515), .ZN(n4488)
         );
  OAI21_X1 U5595 ( .B1(n4844), .B2(n4517), .A(n4488), .ZN(n4489) );
  AOI21_X1 U5596 ( .B1(n6331), .B2(n4519), .A(n4489), .ZN(n4490) );
  OAI21_X1 U5597 ( .B1(n4522), .B2(n4491), .A(n4490), .ZN(U3079) );
  INV_X1 U5598 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4495) );
  AOI22_X1 U5599 ( .A1(n4620), .A2(n6211), .B1(n6360), .B2(n4515), .ZN(n4492)
         );
  OAI21_X1 U5600 ( .B1(n4868), .B2(n4517), .A(n4492), .ZN(n4493) );
  AOI21_X1 U5601 ( .B1(n6356), .B2(n4519), .A(n4493), .ZN(n4494) );
  OAI21_X1 U5602 ( .B1(n4522), .B2(n4495), .A(n4494), .ZN(U3083) );
  INV_X1 U5603 ( .A(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4499) );
  AOI22_X1 U5604 ( .A1(n4620), .A2(n6286), .B1(n6351), .B2(n4515), .ZN(n4496)
         );
  OAI21_X1 U5605 ( .B1(n4856), .B2(n4517), .A(n4496), .ZN(n4497) );
  AOI21_X1 U5606 ( .B1(n6349), .B2(n4519), .A(n4497), .ZN(n4498) );
  OAI21_X1 U5607 ( .B1(n4522), .B2(n4499), .A(n4498), .ZN(U3082) );
  INV_X1 U5608 ( .A(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4503) );
  AOI22_X1 U5609 ( .A1(n4620), .A2(n6282), .B1(n6345), .B2(n4515), .ZN(n4500)
         );
  OAI21_X1 U5610 ( .B1(n4852), .B2(n4517), .A(n4500), .ZN(n4501) );
  AOI21_X1 U5611 ( .B1(n6343), .B2(n4519), .A(n4501), .ZN(n4502) );
  OAI21_X1 U5612 ( .B1(n4522), .B2(n4503), .A(n4502), .ZN(U3081) );
  AOI22_X1 U5613 ( .A1(n4620), .A2(n6270), .B1(n6327), .B2(n4515), .ZN(n4504)
         );
  OAI21_X1 U5614 ( .B1(n4848), .B2(n4517), .A(n4504), .ZN(n4505) );
  AOI21_X1 U5615 ( .B1(n6325), .B2(n4519), .A(n4505), .ZN(n4506) );
  OAI21_X1 U5616 ( .B1(n4522), .B2(n6584), .A(n4506), .ZN(U3078) );
  INV_X1 U5617 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4510) );
  AOI22_X1 U5618 ( .A1(n4620), .A2(n6266), .B1(n6321), .B2(n4515), .ZN(n4507)
         );
  OAI21_X1 U5619 ( .B1(n4860), .B2(n4517), .A(n4507), .ZN(n4508) );
  AOI21_X1 U5620 ( .B1(n6319), .B2(n4519), .A(n4508), .ZN(n4509) );
  OAI21_X1 U5621 ( .B1(n4522), .B2(n4510), .A(n4509), .ZN(U3077) );
  INV_X1 U5622 ( .A(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4514) );
  AOI22_X1 U5623 ( .A1(n4620), .A2(n6185), .B1(n6315), .B2(n4515), .ZN(n4511)
         );
  OAI21_X1 U5624 ( .B1(n4864), .B2(n4517), .A(n4511), .ZN(n4512) );
  AOI21_X1 U5625 ( .B1(n6303), .B2(n4519), .A(n4512), .ZN(n4513) );
  OAI21_X1 U5626 ( .B1(n4522), .B2(n4514), .A(n4513), .ZN(U3076) );
  INV_X1 U5627 ( .A(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4521) );
  AOI22_X1 U5628 ( .A1(n4620), .A2(n6278), .B1(n6339), .B2(n4515), .ZN(n4516)
         );
  OAI21_X1 U5629 ( .B1(n4876), .B2(n4517), .A(n4516), .ZN(n4518) );
  AOI21_X1 U5630 ( .B1(n6337), .B2(n4519), .A(n4518), .ZN(n4520) );
  OAI21_X1 U5631 ( .B1(n4522), .B2(n4521), .A(n4520), .ZN(U3080) );
  NAND3_X1 U5632 ( .A1(n6383), .A2(n6376), .A3(n6372), .ZN(n5706) );
  NOR2_X1 U5633 ( .A1(n4761), .A2(n5706), .ZN(n4524) );
  INV_X1 U5634 ( .A(n4524), .ZN(n4550) );
  NAND2_X1 U5635 ( .A1(n4894), .A2(n5693), .ZN(n5751) );
  OR2_X1 U5636 ( .A1(n4523), .A2(n5751), .ZN(n5704) );
  INV_X1 U5637 ( .A(n5704), .ZN(n5713) );
  AOI21_X1 U5638 ( .B1(n5713), .B2(n6256), .A(n4524), .ZN(n4530) );
  NAND3_X1 U5639 ( .A1(n6188), .A2(n6187), .A3(n4525), .ZN(n4531) );
  OR2_X1 U5640 ( .A1(n4531), .A2(n6305), .ZN(n4526) );
  AND2_X1 U5641 ( .A1(n4526), .A2(n6500), .ZN(n4528) );
  AOI22_X1 U5642 ( .A1(n4530), .A2(n4528), .B1(n6308), .B2(n5706), .ZN(n4527)
         );
  NAND2_X1 U5643 ( .A1(n6259), .A2(n4527), .ZN(n4547) );
  INV_X1 U5644 ( .A(n4528), .ZN(n4529) );
  OAI22_X1 U5645 ( .A1(n4530), .A2(n4529), .B1(n6405), .B2(n5706), .ZN(n4546)
         );
  AOI22_X1 U5646 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4547), .B1(n6343), 
        .B2(n4546), .ZN(n4533) );
  NOR2_X2 U5647 ( .A1(n4531), .A2(n4766), .ZN(n5745) );
  NOR2_X2 U5648 ( .A1(n4531), .A2(n4615), .ZN(n4873) );
  AOI22_X1 U5649 ( .A1(n6282), .A2(n5745), .B1(n4873), .B2(n6345), .ZN(n4532)
         );
  OAI211_X1 U5650 ( .C1(n4852), .C2(n4550), .A(n4533), .B(n4532), .ZN(U3033)
         );
  AOI22_X1 U5651 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4547), .B1(n6337), 
        .B2(n4546), .ZN(n4535) );
  AOI22_X1 U5652 ( .A1(n6278), .A2(n5745), .B1(n4873), .B2(n6339), .ZN(n4534)
         );
  OAI211_X1 U5653 ( .C1(n4876), .C2(n4550), .A(n4535), .B(n4534), .ZN(U3032)
         );
  AOI22_X1 U5654 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4547), .B1(n6325), 
        .B2(n4546), .ZN(n4537) );
  AOI22_X1 U5655 ( .A1(n6270), .A2(n5745), .B1(n4873), .B2(n6327), .ZN(n4536)
         );
  OAI211_X1 U5656 ( .C1(n4848), .C2(n4550), .A(n4537), .B(n4536), .ZN(U3030)
         );
  AOI22_X1 U5657 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4547), .B1(n6349), 
        .B2(n4546), .ZN(n4539) );
  AOI22_X1 U5658 ( .A1(n6286), .A2(n5745), .B1(n4873), .B2(n6351), .ZN(n4538)
         );
  OAI211_X1 U5659 ( .C1(n4856), .C2(n4550), .A(n4539), .B(n4538), .ZN(U3034)
         );
  AOI22_X1 U5660 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4547), .B1(n6356), 
        .B2(n4546), .ZN(n4541) );
  AOI22_X1 U5661 ( .A1(n6211), .A2(n5745), .B1(n4873), .B2(n6360), .ZN(n4540)
         );
  OAI211_X1 U5662 ( .C1(n4868), .C2(n4550), .A(n4541), .B(n4540), .ZN(U3035)
         );
  AOI22_X1 U5663 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4547), .B1(n6303), 
        .B2(n4546), .ZN(n4543) );
  AOI22_X1 U5664 ( .A1(n6185), .A2(n5745), .B1(n4873), .B2(n6315), .ZN(n4542)
         );
  OAI211_X1 U5665 ( .C1(n4864), .C2(n4550), .A(n4543), .B(n4542), .ZN(U3028)
         );
  AOI22_X1 U5666 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4547), .B1(n6319), 
        .B2(n4546), .ZN(n4545) );
  AOI22_X1 U5667 ( .A1(n6266), .A2(n5745), .B1(n4873), .B2(n6321), .ZN(n4544)
         );
  OAI211_X1 U5668 ( .C1(n4860), .C2(n4550), .A(n4545), .B(n4544), .ZN(U3029)
         );
  AOI22_X1 U5669 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4547), .B1(n6331), 
        .B2(n4546), .ZN(n4549) );
  AOI22_X1 U5670 ( .A1(n6274), .A2(n5745), .B1(n4873), .B2(n6333), .ZN(n4548)
         );
  OAI211_X1 U5671 ( .C1(n4844), .C2(n4550), .A(n4549), .B(n4548), .ZN(U3031)
         );
  NAND3_X1 U5672 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6376), .A3(n6372), .ZN(n5754) );
  NOR2_X1 U5673 ( .A1(n4761), .A2(n5754), .ZN(n4551) );
  INV_X1 U5674 ( .A(n4551), .ZN(n4580) );
  INV_X1 U5675 ( .A(n5751), .ZN(n4552) );
  AOI21_X1 U5676 ( .B1(n4553), .B2(n4552), .A(n4551), .ZN(n4558) );
  AOI21_X1 U5677 ( .B1(n4560), .B2(STATEBS16_REG_SCAN_IN), .A(n6308), .ZN(
        n4556) );
  AOI22_X1 U5678 ( .A1(n4558), .A2(n4556), .B1(n6308), .B2(n5754), .ZN(n4555)
         );
  NAND2_X1 U5679 ( .A1(n6259), .A2(n4555), .ZN(n4576) );
  INV_X1 U5680 ( .A(n4556), .ZN(n4557) );
  OAI22_X1 U5681 ( .A1(n4558), .A2(n4557), .B1(n6405), .B2(n5754), .ZN(n4575)
         );
  AOI22_X1 U5682 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4576), .B1(n6303), 
        .B2(n4575), .ZN(n4562) );
  INV_X1 U5683 ( .A(n4560), .ZN(n4559) );
  NAND2_X1 U5684 ( .A1(n4560), .A2(n4766), .ZN(n4754) );
  AOI22_X1 U5685 ( .A1(n5764), .A2(n6185), .B1(n4577), .B2(n6315), .ZN(n4561)
         );
  OAI211_X1 U5686 ( .C1(n4864), .C2(n4580), .A(n4562), .B(n4561), .ZN(U3092)
         );
  AOI22_X1 U5687 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4576), .B1(n6356), 
        .B2(n4575), .ZN(n4564) );
  AOI22_X1 U5688 ( .A1(n5764), .A2(n6211), .B1(n4577), .B2(n6360), .ZN(n4563)
         );
  OAI211_X1 U5689 ( .C1(n4868), .C2(n4580), .A(n4564), .B(n4563), .ZN(U3099)
         );
  AOI22_X1 U5690 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4576), .B1(n6349), 
        .B2(n4575), .ZN(n4566) );
  AOI22_X1 U5691 ( .A1(n5764), .A2(n6286), .B1(n4577), .B2(n6351), .ZN(n4565)
         );
  OAI211_X1 U5692 ( .C1(n4856), .C2(n4580), .A(n4566), .B(n4565), .ZN(U3098)
         );
  AOI22_X1 U5693 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4576), .B1(n6343), 
        .B2(n4575), .ZN(n4568) );
  AOI22_X1 U5694 ( .A1(n5764), .A2(n6282), .B1(n4577), .B2(n6345), .ZN(n4567)
         );
  OAI211_X1 U5695 ( .C1(n4852), .C2(n4580), .A(n4568), .B(n4567), .ZN(U3097)
         );
  AOI22_X1 U5696 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4576), .B1(n6337), 
        .B2(n4575), .ZN(n4570) );
  AOI22_X1 U5697 ( .A1(n5764), .A2(n6278), .B1(n4577), .B2(n6339), .ZN(n4569)
         );
  OAI211_X1 U5698 ( .C1(n4876), .C2(n4580), .A(n4570), .B(n4569), .ZN(U3096)
         );
  AOI22_X1 U5699 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4576), .B1(n6331), 
        .B2(n4575), .ZN(n4572) );
  AOI22_X1 U5700 ( .A1(n5764), .A2(n6274), .B1(n4577), .B2(n6333), .ZN(n4571)
         );
  OAI211_X1 U5701 ( .C1(n4844), .C2(n4580), .A(n4572), .B(n4571), .ZN(U3095)
         );
  AOI22_X1 U5702 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4576), .B1(n6319), 
        .B2(n4575), .ZN(n4574) );
  AOI22_X1 U5703 ( .A1(n5764), .A2(n6266), .B1(n4577), .B2(n6321), .ZN(n4573)
         );
  OAI211_X1 U5704 ( .C1(n4860), .C2(n4580), .A(n4574), .B(n4573), .ZN(U3093)
         );
  AOI22_X1 U5705 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4576), .B1(n6325), 
        .B2(n4575), .ZN(n4579) );
  AOI22_X1 U5706 ( .A1(n5764), .A2(n6270), .B1(n4577), .B2(n6327), .ZN(n4578)
         );
  OAI211_X1 U5707 ( .C1(n4848), .C2(n4580), .A(n4579), .B(n4578), .ZN(U3094)
         );
  OAI21_X1 U5708 ( .B1(n4582), .B2(n4581), .A(n4719), .ZN(n4714) );
  AOI22_X1 U5709 ( .A1(n5544), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n6014), .ZN(n4583) );
  OAI21_X1 U5710 ( .B1(n4714), .B2(n5862), .A(n4583), .ZN(U2883) );
  INV_X1 U5711 ( .A(n4914), .ZN(n4587) );
  OAI21_X1 U5712 ( .B1(n5978), .B2(n4587), .A(n4992), .ZN(n5960) );
  NAND2_X1 U5713 ( .A1(n4671), .A2(n4584), .ZN(n4878) );
  OAI21_X1 U5714 ( .B1(n4584), .B2(n4671), .A(n4878), .ZN(n4700) );
  INV_X1 U5715 ( .A(n4585), .ZN(n4586) );
  NOR3_X1 U5716 ( .A1(n5978), .A2(n4587), .A3(n4586), .ZN(n4588) );
  AOI21_X1 U5717 ( .B1(EBX_REG_8__SCAN_IN), .B2(n5993), .A(n4588), .ZN(n4590)
         );
  INV_X1 U5718 ( .A(n5982), .ZN(n5956) );
  AOI21_X1 U5719 ( .B1(n5991), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n5956), 
        .ZN(n4589) );
  OAI211_X1 U5720 ( .C1(n5983), .C2(n4700), .A(n4590), .B(n4589), .ZN(n4591)
         );
  AOI21_X1 U5721 ( .B1(REIP_REG_8__SCAN_IN), .B2(n5960), .A(n4591), .ZN(n4593)
         );
  NAND2_X1 U5722 ( .A1(n5958), .A2(n4713), .ZN(n4592) );
  OAI211_X1 U5723 ( .C1(n4714), .C2(n5820), .A(n4593), .B(n4592), .ZN(U2819)
         );
  INV_X1 U5724 ( .A(n4594), .ZN(n4596) );
  XNOR2_X1 U5725 ( .A(n4596), .B(n4595), .ZN(n6089) );
  INV_X1 U5726 ( .A(n6089), .ZN(n4675) );
  INV_X1 U5727 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6029) );
  OAI222_X1 U5728 ( .A1(n5862), .A2(n4675), .B1(n5127), .B2(n4597), .C1(n5421), 
        .C2(n6029), .ZN(U2884) );
  INV_X1 U5729 ( .A(n4602), .ZN(n4598) );
  OAI21_X1 U5730 ( .B1(n4599), .B2(n4598), .A(n5820), .ZN(n6000) );
  INV_X1 U5731 ( .A(n6000), .ZN(n4902) );
  INV_X1 U5732 ( .A(n4600), .ZN(n4601) );
  NAND2_X1 U5733 ( .A1(n4602), .A2(n4601), .ZN(n5996) );
  INV_X1 U5734 ( .A(n4603), .ZN(n6154) );
  OAI21_X1 U5735 ( .B1(n4890), .B2(n4605), .A(n5459), .ZN(n6003) );
  OAI22_X1 U5736 ( .A1(n6003), .A2(n6436), .B1(n4663), .B2(n5815), .ZN(n4604)
         );
  AOI211_X1 U5737 ( .C1(n5992), .C2(n6154), .A(n4604), .B(n5956), .ZN(n4608)
         );
  NOR3_X1 U5738 ( .A1(n5978), .A2(REIP_REG_4__SCAN_IN), .A3(n4605), .ZN(n4606)
         );
  AOI21_X1 U5739 ( .B1(n5993), .B2(EBX_REG_4__SCAN_IN), .A(n4606), .ZN(n4607)
         );
  OAI211_X1 U5740 ( .C1(n4609), .C2(n5996), .A(n4608), .B(n4607), .ZN(n4610)
         );
  AOI21_X1 U5741 ( .B1(n5958), .B2(n4667), .A(n4610), .ZN(n4611) );
  OAI21_X1 U5742 ( .B1(n4902), .B2(n4664), .A(n4611), .ZN(U2823) );
  NAND2_X1 U5743 ( .A1(n4761), .A2(n4612), .ZN(n4652) );
  NOR2_X1 U5744 ( .A1(n4554), .A2(n5696), .ZN(n4613) );
  NAND2_X1 U5745 ( .A1(n4614), .A2(n4613), .ZN(n4767) );
  NOR3_X1 U5746 ( .A1(n4649), .A2(n4620), .A3(n6308), .ZN(n4616) );
  OAI21_X1 U5747 ( .B1(n4616), .B2(n6224), .A(n4621), .ZN(n4619) );
  AOI21_X1 U5748 ( .B1(n4652), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4617) );
  NAND3_X1 U5749 ( .A1(n4619), .A2(n4618), .A3(n4617), .ZN(n4645) );
  NAND2_X1 U5750 ( .A1(n4645), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4626) );
  INV_X1 U5751 ( .A(n4620), .ZN(n4647) );
  NOR2_X1 U5752 ( .A1(n6300), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4623)
         );
  NOR3_X1 U5753 ( .A1(n6222), .A2(n4621), .A3(n6308), .ZN(n4622) );
  AOI21_X1 U5754 ( .B1(n5756), .B2(n4623), .A(n4622), .ZN(n4646) );
  OAI22_X1 U5755 ( .A1(n4647), .A2(n6285), .B1(n4646), .B2(n5788), .ZN(n4624)
         );
  AOI21_X1 U5756 ( .B1(n6282), .B2(n4649), .A(n4624), .ZN(n4625) );
  OAI211_X1 U5757 ( .C1(n4652), .C2(n4852), .A(n4626), .B(n4625), .ZN(U3073)
         );
  NAND2_X1 U5758 ( .A1(n4645), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4629) );
  OAI22_X1 U5759 ( .A1(n4647), .A2(n6218), .B1(n4646), .B2(n5798), .ZN(n4627)
         );
  AOI21_X1 U5760 ( .B1(n6211), .B2(n4649), .A(n4627), .ZN(n4628) );
  OAI211_X1 U5761 ( .C1(n4652), .C2(n4868), .A(n4629), .B(n4628), .ZN(U3075)
         );
  NAND2_X1 U5762 ( .A1(n4645), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4632) );
  OAI22_X1 U5763 ( .A1(n4647), .A2(n6269), .B1(n4646), .B2(n5768), .ZN(n4630)
         );
  AOI21_X1 U5764 ( .B1(n6266), .B2(n4649), .A(n4630), .ZN(n4631) );
  OAI211_X1 U5765 ( .C1(n4652), .C2(n4860), .A(n4632), .B(n4631), .ZN(U3069)
         );
  NAND2_X1 U5766 ( .A1(n4645), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4635) );
  OAI22_X1 U5767 ( .A1(n4647), .A2(n6277), .B1(n4646), .B2(n5778), .ZN(n4633)
         );
  AOI21_X1 U5768 ( .B1(n6274), .B2(n4649), .A(n4633), .ZN(n4634) );
  OAI211_X1 U5769 ( .C1(n4652), .C2(n4844), .A(n4635), .B(n4634), .ZN(U3071)
         );
  NAND2_X1 U5770 ( .A1(n4645), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4638) );
  OAI22_X1 U5771 ( .A1(n4647), .A2(n6290), .B1(n4646), .B2(n5793), .ZN(n4636)
         );
  AOI21_X1 U5772 ( .B1(n6286), .B2(n4649), .A(n4636), .ZN(n4637) );
  OAI211_X1 U5773 ( .C1(n4652), .C2(n4856), .A(n4638), .B(n4637), .ZN(U3074)
         );
  NAND2_X1 U5774 ( .A1(n4645), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4641) );
  OAI22_X1 U5775 ( .A1(n4647), .A2(n6281), .B1(n4646), .B2(n5783), .ZN(n4639)
         );
  AOI21_X1 U5776 ( .B1(n6278), .B2(n4649), .A(n4639), .ZN(n4640) );
  OAI211_X1 U5777 ( .C1(n4652), .C2(n4876), .A(n4641), .B(n4640), .ZN(U3072)
         );
  NAND2_X1 U5778 ( .A1(n4645), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4644) );
  OAI22_X1 U5779 ( .A1(n4647), .A2(n6198), .B1(n4646), .B2(n5762), .ZN(n4642)
         );
  AOI21_X1 U5780 ( .B1(n6185), .B2(n4649), .A(n4642), .ZN(n4643) );
  OAI211_X1 U5781 ( .C1(n4864), .C2(n4652), .A(n4644), .B(n4643), .ZN(U3068)
         );
  NAND2_X1 U5782 ( .A1(n4645), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4651) );
  OAI22_X1 U5783 ( .A1(n4647), .A2(n6273), .B1(n4646), .B2(n5773), .ZN(n4648)
         );
  AOI21_X1 U5784 ( .B1(n6270), .B2(n4649), .A(n4648), .ZN(n4650) );
  OAI211_X1 U5785 ( .C1(n4652), .C2(n4848), .A(n4651), .B(n4650), .ZN(U3070)
         );
  AND2_X1 U5786 ( .A1(n5993), .A2(EBX_REG_0__SCAN_IN), .ZN(n4656) );
  OAI22_X1 U5787 ( .A1(n4654), .A2(n5996), .B1(n5983), .B2(n4653), .ZN(n4655)
         );
  AOI211_X1 U5788 ( .C1(REIP_REG_0__SCAN_IN), .C2(n5459), .A(n4656), .B(n4655), 
        .ZN(n4658) );
  OAI21_X1 U5789 ( .B1(n5958), .B2(n5991), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4657) );
  OAI211_X1 U5790 ( .C1(n4902), .C2(n4659), .A(n4658), .B(n4657), .ZN(U2827)
         );
  OAI21_X1 U5791 ( .B1(n4662), .B2(n4661), .A(n4660), .ZN(n6152) );
  OAI22_X1 U5792 ( .A1(n5597), .A2(n4663), .B1(n5585), .B2(n6436), .ZN(n4666)
         );
  NOR2_X1 U5793 ( .A1(n4664), .A2(n5591), .ZN(n4665) );
  AOI211_X1 U5794 ( .C1(n5593), .C2(n4667), .A(n4666), .B(n4665), .ZN(n4668)
         );
  OAI21_X1 U5795 ( .B1(n5912), .B2(n6152), .A(n4668), .ZN(U2982) );
  OAI222_X1 U5796 ( .A1(n4700), .A2(n5535), .B1(n5532), .B2(n3043), .C1(n2945), 
        .C2(n4714), .ZN(U2851) );
  NAND2_X1 U5797 ( .A1(n4670), .A2(n4669), .ZN(n4673) );
  INV_X1 U5798 ( .A(n4671), .ZN(n4672) );
  NAND2_X1 U5799 ( .A1(n4673), .A2(n4672), .ZN(n6135) );
  INV_X1 U5800 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4674) );
  OAI222_X1 U5801 ( .A1(n6135), .A2(n5535), .B1(n2945), .B2(n4675), .C1(n5532), 
        .C2(n4674), .ZN(U2852) );
  NAND2_X1 U5802 ( .A1(n4677), .A2(n4676), .ZN(n4683) );
  INV_X1 U5803 ( .A(n4678), .ZN(n4680) );
  NAND2_X1 U5804 ( .A1(n4680), .A2(n4679), .ZN(n4695) );
  XNOR2_X1 U5805 ( .A(n4695), .B(n4696), .ZN(n4681) );
  NAND2_X1 U5806 ( .A1(n4681), .A2(n4697), .ZN(n4682) );
  INV_X1 U5807 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6141) );
  XNOR2_X1 U5808 ( .A(n4689), .B(n6141), .ZN(n6086) );
  AND2_X1 U5809 ( .A1(n4684), .A2(n6086), .ZN(n4687) );
  XNOR2_X1 U5810 ( .A(n4689), .B(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4686)
         );
  NAND2_X1 U5811 ( .A1(n4685), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6083)
         );
  AOI21_X2 U5812 ( .B1(n4688), .B2(n4687), .A(n2952), .ZN(n6085) );
  NAND2_X1 U5813 ( .A1(n4689), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4690)
         );
  NAND2_X1 U5814 ( .A1(n6085), .A2(n4690), .ZN(n4803) );
  NOR2_X1 U5815 ( .A1(n4692), .A2(n4691), .ZN(n4693) );
  NAND2_X4 U5816 ( .A1(n4694), .A2(n4693), .ZN(n5581) );
  INV_X1 U5817 ( .A(n4695), .ZN(n4698) );
  NAND3_X1 U5818 ( .A1(n4698), .A2(n4697), .A3(n4696), .ZN(n4699) );
  INV_X1 U5819 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4705) );
  XNOR2_X1 U5820 ( .A(n4805), .B(n4705), .ZN(n4800) );
  NAND2_X1 U5821 ( .A1(n5001), .A2(n4800), .ZN(n4926) );
  OAI21_X1 U5822 ( .B1(n5001), .B2(n4800), .A(n4926), .ZN(n4718) );
  INV_X1 U5823 ( .A(n4700), .ZN(n4708) );
  INV_X1 U5824 ( .A(REIP_REG_8__SCAN_IN), .ZN(n4701) );
  NOR2_X1 U5825 ( .A1(n5585), .A2(n4701), .ZN(n4712) );
  NOR2_X1 U5826 ( .A1(n6141), .A2(n4705), .ZN(n4934) );
  NAND3_X1 U5827 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6144), .ZN(n4816) );
  NOR2_X1 U5828 ( .A1(n6155), .A2(n4816), .ZN(n6137) );
  OAI21_X1 U5829 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6137), .ZN(n4706) );
  INV_X1 U5830 ( .A(n6156), .ZN(n4702) );
  NAND4_X1 U5831 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6176), .A4(n4702), .ZN(n4815) );
  INV_X1 U5832 ( .A(n4816), .ZN(n4703) );
  OAI21_X1 U5833 ( .B1(n4703), .B2(n5074), .A(n5054), .ZN(n4704) );
  AOI21_X1 U5834 ( .B1(n5052), .B2(n4815), .A(n4704), .ZN(n6142) );
  OAI22_X1 U5835 ( .A1(n4934), .A2(n4706), .B1(n6142), .B2(n4705), .ZN(n4707)
         );
  AOI211_X1 U5836 ( .C1(n6168), .C2(n4708), .A(n4712), .B(n4707), .ZN(n4709)
         );
  OAI21_X1 U5837 ( .B1(n5680), .B2(n4718), .A(n4709), .ZN(U3010) );
  INV_X1 U5838 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4710) );
  NOR2_X1 U5839 ( .A1(n5597), .A2(n4710), .ZN(n4711) );
  AOI211_X1 U5840 ( .C1(n5593), .C2(n4713), .A(n4712), .B(n4711), .ZN(n4717)
         );
  INV_X1 U5841 ( .A(n4714), .ZN(n4715) );
  NAND2_X1 U5842 ( .A1(n4715), .A2(n2946), .ZN(n4716) );
  OAI211_X1 U5843 ( .C1(n4718), .C2(n5912), .A(n4717), .B(n4716), .ZN(U2978)
         );
  INV_X1 U5844 ( .A(n4719), .ZN(n4723) );
  INV_X1 U5845 ( .A(n4720), .ZN(n4722) );
  OAI21_X1 U5846 ( .B1(n4723), .B2(n4722), .A(n4921), .ZN(n4911) );
  AOI22_X1 U5847 ( .A1(n5544), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n6014), .ZN(n4724) );
  OAI21_X1 U5848 ( .B1(n4911), .B2(n5862), .A(n4724), .ZN(U2882) );
  AOI21_X1 U5849 ( .B1(n4754), .B2(n6297), .A(n6305), .ZN(n4725) );
  NOR2_X1 U5850 ( .A1(n4725), .A2(n6308), .ZN(n4730) );
  AND2_X1 U5851 ( .A1(n4894), .A2(n4886), .ZN(n4834) );
  AND2_X1 U5852 ( .A1(n4834), .A2(n6222), .ZN(n6257) );
  INV_X1 U5853 ( .A(n6226), .ZN(n6312) );
  NOR2_X1 U5854 ( .A1(n6312), .A2(n6383), .ZN(n4726) );
  AOI22_X1 U5855 ( .A1(n4730), .A2(n6257), .B1(n5756), .B2(n4726), .ZN(n4759)
         );
  NAND3_X1 U5856 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6376), .ZN(n6261) );
  NOR2_X1 U5857 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6261), .ZN(n4756)
         );
  NOR2_X1 U5858 ( .A1(n5709), .A2(n4727), .ZN(n4837) );
  INV_X1 U5859 ( .A(n6257), .ZN(n4729) );
  AOI21_X1 U5860 ( .B1(n4730), .B2(n4729), .A(n4728), .ZN(n4731) );
  OAI211_X1 U5861 ( .C1(n4756), .C2(n6483), .A(n4837), .B(n4731), .ZN(n4753)
         );
  NAND2_X1 U5862 ( .A1(n4753), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4734)
         );
  OAI22_X1 U5863 ( .A1(n4754), .A2(n6324), .B1(n6297), .B2(n6269), .ZN(n4732)
         );
  AOI21_X1 U5864 ( .B1(n4756), .B2(n6320), .A(n4732), .ZN(n4733) );
  OAI211_X1 U5865 ( .C1(n4759), .C2(n5768), .A(n4734), .B(n4733), .ZN(U3101)
         );
  NAND2_X1 U5866 ( .A1(n4753), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4737)
         );
  OAI22_X1 U5867 ( .A1(n4754), .A2(n6336), .B1(n6297), .B2(n6277), .ZN(n4735)
         );
  AOI21_X1 U5868 ( .B1(n4756), .B2(n6332), .A(n4735), .ZN(n4736) );
  OAI211_X1 U5869 ( .C1(n4759), .C2(n5778), .A(n4737), .B(n4736), .ZN(U3103)
         );
  NAND2_X1 U5870 ( .A1(n4753), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4740)
         );
  OAI22_X1 U5871 ( .A1(n4754), .A2(n6354), .B1(n6297), .B2(n6290), .ZN(n4738)
         );
  AOI21_X1 U5872 ( .B1(n4756), .B2(n6350), .A(n4738), .ZN(n4739) );
  OAI211_X1 U5873 ( .C1(n4759), .C2(n5793), .A(n4740), .B(n4739), .ZN(U3106)
         );
  NAND2_X1 U5874 ( .A1(n4753), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4743)
         );
  OAI22_X1 U5875 ( .A1(n4754), .A2(n6365), .B1(n6297), .B2(n6218), .ZN(n4741)
         );
  AOI21_X1 U5876 ( .B1(n4756), .B2(n6358), .A(n4741), .ZN(n4742) );
  OAI211_X1 U5877 ( .C1(n4759), .C2(n5798), .A(n4743), .B(n4742), .ZN(U3107)
         );
  NAND2_X1 U5878 ( .A1(n4753), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4746)
         );
  OAI22_X1 U5879 ( .A1(n4754), .A2(n6330), .B1(n6297), .B2(n6273), .ZN(n4744)
         );
  AOI21_X1 U5880 ( .B1(n4756), .B2(n6326), .A(n4744), .ZN(n4745) );
  OAI211_X1 U5881 ( .C1(n4759), .C2(n5773), .A(n4746), .B(n4745), .ZN(U3102)
         );
  NAND2_X1 U5882 ( .A1(n4753), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4749)
         );
  OAI22_X1 U5883 ( .A1(n4754), .A2(n6348), .B1(n6297), .B2(n6285), .ZN(n4747)
         );
  AOI21_X1 U5884 ( .B1(n4756), .B2(n6344), .A(n4747), .ZN(n4748) );
  OAI211_X1 U5885 ( .C1(n4759), .C2(n5788), .A(n4749), .B(n4748), .ZN(U3105)
         );
  NAND2_X1 U5886 ( .A1(n4753), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4752)
         );
  OAI22_X1 U5887 ( .A1(n4754), .A2(n6342), .B1(n6297), .B2(n6281), .ZN(n4750)
         );
  AOI21_X1 U5888 ( .B1(n4756), .B2(n6338), .A(n4750), .ZN(n4751) );
  OAI211_X1 U5889 ( .C1(n4759), .C2(n5783), .A(n4752), .B(n4751), .ZN(U3104)
         );
  NAND2_X1 U5890 ( .A1(n4753), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4758)
         );
  OAI22_X1 U5891 ( .A1(n4754), .A2(n6318), .B1(n6297), .B2(n6198), .ZN(n4755)
         );
  AOI21_X1 U5892 ( .B1(n4756), .B2(n6304), .A(n4755), .ZN(n4757) );
  OAI211_X1 U5893 ( .C1(n4759), .C2(n5762), .A(n4758), .B(n4757), .ZN(U3100)
         );
  OAI21_X1 U5894 ( .B1(n4767), .B2(n6305), .A(n6500), .ZN(n6230) );
  INV_X1 U5895 ( .A(n6230), .ZN(n4765) );
  NAND2_X1 U5896 ( .A1(n4760), .A2(n6383), .ZN(n6219) );
  NOR2_X1 U5897 ( .A1(n4761), .A2(n6219), .ZN(n4794) );
  INV_X1 U5898 ( .A(n4794), .ZN(n4762) );
  OAI21_X1 U5899 ( .B1(n6223), .B2(n4763), .A(n4762), .ZN(n4770) );
  INV_X1 U5900 ( .A(n6219), .ZN(n4764) );
  AOI22_X1 U5901 ( .A1(n4765), .A2(n4770), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4764), .ZN(n4798) );
  NOR2_X1 U5902 ( .A1(n4767), .A2(n4766), .ZN(n6247) );
  INV_X1 U5903 ( .A(n6247), .ZN(n4792) );
  OAI22_X1 U5904 ( .A1(n4792), .A2(n6365), .B1(n6218), .B2(n4791), .ZN(n4768)
         );
  AOI21_X1 U5905 ( .B1(n6358), .B2(n4794), .A(n4768), .ZN(n4772) );
  NAND2_X1 U5906 ( .A1(n6219), .A2(n6308), .ZN(n4769) );
  OAI211_X1 U5907 ( .C1(n6230), .C2(n4770), .A(n6259), .B(n4769), .ZN(n4795)
         );
  NAND2_X1 U5908 ( .A1(n4795), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4771) );
  OAI211_X1 U5909 ( .C1(n4798), .C2(n5798), .A(n4772), .B(n4771), .ZN(U3067)
         );
  OAI22_X1 U5910 ( .A1(n4792), .A2(n6336), .B1(n6277), .B2(n4791), .ZN(n4773)
         );
  AOI21_X1 U5911 ( .B1(n6332), .B2(n4794), .A(n4773), .ZN(n4775) );
  NAND2_X1 U5912 ( .A1(n4795), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4774) );
  OAI211_X1 U5913 ( .C1(n4798), .C2(n5778), .A(n4775), .B(n4774), .ZN(U3063)
         );
  OAI22_X1 U5914 ( .A1(n4792), .A2(n6318), .B1(n6198), .B2(n4791), .ZN(n4776)
         );
  AOI21_X1 U5915 ( .B1(n6304), .B2(n4794), .A(n4776), .ZN(n4778) );
  NAND2_X1 U5916 ( .A1(n4795), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4777) );
  OAI211_X1 U5917 ( .C1(n4798), .C2(n5762), .A(n4778), .B(n4777), .ZN(U3060)
         );
  OAI22_X1 U5918 ( .A1(n4792), .A2(n6324), .B1(n6269), .B2(n4791), .ZN(n4779)
         );
  AOI21_X1 U5919 ( .B1(n6320), .B2(n4794), .A(n4779), .ZN(n4781) );
  NAND2_X1 U5920 ( .A1(n4795), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4780) );
  OAI211_X1 U5921 ( .C1(n4798), .C2(n5768), .A(n4781), .B(n4780), .ZN(U3061)
         );
  OAI22_X1 U5922 ( .A1(n4792), .A2(n6330), .B1(n6273), .B2(n4791), .ZN(n4782)
         );
  AOI21_X1 U5923 ( .B1(n6326), .B2(n4794), .A(n4782), .ZN(n4784) );
  NAND2_X1 U5924 ( .A1(n4795), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4783) );
  OAI211_X1 U5925 ( .C1(n4798), .C2(n5773), .A(n4784), .B(n4783), .ZN(U3062)
         );
  OAI22_X1 U5926 ( .A1(n4792), .A2(n6348), .B1(n6285), .B2(n4791), .ZN(n4785)
         );
  AOI21_X1 U5927 ( .B1(n6344), .B2(n4794), .A(n4785), .ZN(n4787) );
  NAND2_X1 U5928 ( .A1(n4795), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4786) );
  OAI211_X1 U5929 ( .C1(n4798), .C2(n5788), .A(n4787), .B(n4786), .ZN(U3065)
         );
  OAI22_X1 U5930 ( .A1(n4792), .A2(n6342), .B1(n6281), .B2(n4791), .ZN(n4788)
         );
  AOI21_X1 U5931 ( .B1(n6338), .B2(n4794), .A(n4788), .ZN(n4790) );
  NAND2_X1 U5932 ( .A1(n4795), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4789) );
  OAI211_X1 U5933 ( .C1(n4798), .C2(n5783), .A(n4790), .B(n4789), .ZN(U3064)
         );
  OAI22_X1 U5934 ( .A1(n4792), .A2(n6354), .B1(n6290), .B2(n4791), .ZN(n4793)
         );
  AOI21_X1 U5935 ( .B1(n6350), .B2(n4794), .A(n4793), .ZN(n4797) );
  NAND2_X1 U5936 ( .A1(n4795), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4796) );
  OAI211_X1 U5937 ( .C1(n4798), .C2(n5793), .A(n4797), .B(n4796), .ZN(U3066)
         );
  INV_X1 U5938 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4799) );
  NAND2_X1 U5939 ( .A1(n5581), .A2(n4799), .ZN(n4924) );
  INV_X1 U5940 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6515) );
  NAND2_X1 U5941 ( .A1(n5581), .A2(n6515), .ZN(n4927) );
  AND2_X1 U5942 ( .A1(n4924), .A2(n4927), .ZN(n4804) );
  AND2_X1 U5943 ( .A1(n4800), .A2(n4804), .ZN(n5000) );
  INV_X1 U5944 ( .A(n4807), .ZN(n4801) );
  AND2_X1 U5945 ( .A1(n5000), .A2(n4801), .ZN(n4802) );
  NAND2_X1 U5946 ( .A1(n4803), .A2(n4802), .ZN(n4809) );
  INV_X1 U5947 ( .A(n4804), .ZN(n4806) );
  NAND2_X1 U5948 ( .A1(n4805), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4903)
         );
  NAND2_X1 U5949 ( .A1(n4811), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4904)
         );
  AND2_X1 U5950 ( .A1(n4903), .A2(n4904), .ZN(n4925) );
  AND2_X2 U5951 ( .A1(n4809), .A2(n4808), .ZN(n4942) );
  NAND2_X1 U5952 ( .A1(n4811), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5004) );
  NAND2_X1 U5953 ( .A1(n5875), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4810) );
  NAND2_X1 U5954 ( .A1(n4942), .A2(n4940), .ZN(n4814) );
  INV_X1 U5955 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4826) );
  NOR2_X1 U5956 ( .A1(n5581), .A2(n4826), .ZN(n4938) );
  NAND2_X1 U5957 ( .A1(n5581), .A2(n4826), .ZN(n4959) );
  INV_X1 U5958 ( .A(n4959), .ZN(n4812) );
  NOR2_X1 U5959 ( .A1(n4938), .A2(n4812), .ZN(n4813) );
  XNOR2_X1 U5960 ( .A(n4814), .B(n4813), .ZN(n5135) );
  INV_X1 U5961 ( .A(n5054), .ZN(n4820) );
  NAND3_X1 U5962 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n4934), .ZN(n4817) );
  NOR2_X1 U5963 ( .A1(n4815), .A2(n4817), .ZN(n5049) );
  NOR2_X1 U5964 ( .A1(n4817), .A2(n4816), .ZN(n5050) );
  OAI22_X1 U5965 ( .A1(n4818), .A2(n5049), .B1(n5050), .B2(n5074), .ZN(n4819)
         );
  NOR2_X1 U5966 ( .A1(n4820), .A2(n4819), .ZN(n6127) );
  INV_X1 U5967 ( .A(n6127), .ZN(n4829) );
  INV_X1 U5968 ( .A(n6168), .ZN(n5655) );
  AND2_X1 U5969 ( .A1(n4821), .A2(n4931), .ZN(n4985) );
  OAI21_X1 U5970 ( .B1(n4822), .B2(n4985), .A(n5137), .ZN(n5088) );
  NAND2_X1 U5971 ( .A1(n6167), .A2(REIP_REG_12__SCAN_IN), .ZN(n5128) );
  OAI21_X1 U5972 ( .B1(n5655), .B2(n5088), .A(n5128), .ZN(n4828) );
  INV_X1 U5973 ( .A(n5050), .ZN(n4825) );
  NAND3_X1 U5974 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n4823), .A3(n5049), 
        .ZN(n4824) );
  OAI21_X1 U5975 ( .B1(n4825), .B2(n5074), .A(n4824), .ZN(n4969) );
  AOI21_X1 U5976 ( .B1(n4965), .B2(n5049), .A(n4969), .ZN(n5898) );
  NOR2_X1 U5977 ( .A1(n6126), .A2(n4826), .ZN(n4968) );
  AOI211_X1 U5978 ( .C1(n6126), .C2(n4826), .A(n5898), .B(n4968), .ZN(n4827)
         );
  AOI211_X1 U5979 ( .C1(INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n4829), .A(n4828), .B(n4827), .ZN(n4830) );
  OAI21_X1 U5980 ( .B1(n5135), .B2(n5680), .A(n4830), .ZN(U3006) );
  NAND3_X1 U5981 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6383), .A3(n6376), .ZN(n6193) );
  NOR2_X1 U5982 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6193), .ZN(n4839)
         );
  INV_X1 U5983 ( .A(n4839), .ZN(n4877) );
  NOR2_X1 U5984 ( .A1(n4832), .A2(n4831), .ZN(n4833) );
  NAND2_X1 U5985 ( .A1(n4833), .A2(n6187), .ZN(n4871) );
  OAI21_X1 U5986 ( .B1(n4873), .B2(n6212), .A(n5752), .ZN(n4836) );
  AND2_X1 U5987 ( .A1(n6301), .A2(n4834), .ZN(n6190) );
  INV_X1 U5988 ( .A(n6190), .ZN(n4835) );
  NAND2_X1 U5989 ( .A1(n4836), .A2(n4835), .ZN(n4838) );
  OAI221_X1 U5990 ( .B1(n4839), .B2(n6483), .C1(n4839), .C2(n4838), .A(n4837), 
        .ZN(n4869) );
  NAND2_X1 U5991 ( .A1(n4869), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4843) );
  NOR2_X1 U5992 ( .A1(n6312), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4840)
         );
  AOI22_X1 U5993 ( .A1(n6190), .A2(n6500), .B1(n5756), .B2(n4840), .ZN(n4870)
         );
  OAI22_X1 U5994 ( .A1(n4871), .A2(n6277), .B1(n4870), .B2(n5778), .ZN(n4841)
         );
  AOI21_X1 U5995 ( .B1(n4873), .B2(n6274), .A(n4841), .ZN(n4842) );
  OAI211_X1 U5996 ( .C1(n4877), .C2(n4844), .A(n4843), .B(n4842), .ZN(U3039)
         );
  NAND2_X1 U5997 ( .A1(n4869), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4847) );
  OAI22_X1 U5998 ( .A1(n4871), .A2(n6273), .B1(n4870), .B2(n5773), .ZN(n4845)
         );
  AOI21_X1 U5999 ( .B1(n4873), .B2(n6270), .A(n4845), .ZN(n4846) );
  OAI211_X1 U6000 ( .C1(n4877), .C2(n4848), .A(n4847), .B(n4846), .ZN(U3038)
         );
  NAND2_X1 U6001 ( .A1(n4869), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4851) );
  OAI22_X1 U6002 ( .A1(n4871), .A2(n6285), .B1(n4870), .B2(n5788), .ZN(n4849)
         );
  AOI21_X1 U6003 ( .B1(n4873), .B2(n6282), .A(n4849), .ZN(n4850) );
  OAI211_X1 U6004 ( .C1(n4877), .C2(n4852), .A(n4851), .B(n4850), .ZN(U3041)
         );
  NAND2_X1 U6005 ( .A1(n4869), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4855) );
  OAI22_X1 U6006 ( .A1(n4871), .A2(n6290), .B1(n4870), .B2(n5793), .ZN(n4853)
         );
  AOI21_X1 U6007 ( .B1(n4873), .B2(n6286), .A(n4853), .ZN(n4854) );
  OAI211_X1 U6008 ( .C1(n4877), .C2(n4856), .A(n4855), .B(n4854), .ZN(U3042)
         );
  NAND2_X1 U6009 ( .A1(n4869), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4859) );
  OAI22_X1 U6010 ( .A1(n4871), .A2(n6269), .B1(n4870), .B2(n5768), .ZN(n4857)
         );
  AOI21_X1 U6011 ( .B1(n4873), .B2(n6266), .A(n4857), .ZN(n4858) );
  OAI211_X1 U6012 ( .C1(n4877), .C2(n4860), .A(n4859), .B(n4858), .ZN(U3037)
         );
  NAND2_X1 U6013 ( .A1(n4869), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4863) );
  OAI22_X1 U6014 ( .A1(n4871), .A2(n6198), .B1(n4870), .B2(n5762), .ZN(n4861)
         );
  AOI21_X1 U6015 ( .B1(n4873), .B2(n6185), .A(n4861), .ZN(n4862) );
  OAI211_X1 U6016 ( .C1(n4864), .C2(n4877), .A(n4863), .B(n4862), .ZN(U3036)
         );
  NAND2_X1 U6017 ( .A1(n4869), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4867) );
  OAI22_X1 U6018 ( .A1(n4871), .A2(n6218), .B1(n4870), .B2(n5798), .ZN(n4865)
         );
  AOI21_X1 U6019 ( .B1(n4873), .B2(n6211), .A(n4865), .ZN(n4866) );
  OAI211_X1 U6020 ( .C1(n4877), .C2(n4868), .A(n4867), .B(n4866), .ZN(U3043)
         );
  NAND2_X1 U6021 ( .A1(n4869), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4875) );
  OAI22_X1 U6022 ( .A1(n4871), .A2(n6281), .B1(n4870), .B2(n5783), .ZN(n4872)
         );
  AOI21_X1 U6023 ( .B1(n4873), .B2(n6278), .A(n4872), .ZN(n4874) );
  OAI211_X1 U6024 ( .C1(n4877), .C2(n4876), .A(n4875), .B(n4874), .ZN(U3040)
         );
  NOR2_X1 U6025 ( .A1(n4879), .A2(n4878), .ZN(n4932) );
  AOI21_X1 U6026 ( .B1(n4879), .B2(n4878), .A(n4932), .ZN(n6129) );
  INV_X1 U6027 ( .A(n6129), .ZN(n4881) );
  OAI222_X1 U6028 ( .A1(n4881), .A2(n5535), .B1(n4880), .B2(n5532), .C1(n2945), 
        .C2(n4911), .ZN(U2850) );
  INV_X1 U6029 ( .A(n5996), .ZN(n4887) );
  NOR2_X1 U6030 ( .A1(n5978), .A2(REIP_REG_1__SCAN_IN), .ZN(n4891) );
  AOI21_X1 U6031 ( .B1(EBX_REG_1__SCAN_IN), .B2(n5993), .A(n4891), .ZN(n4883)
         );
  AOI22_X1 U6032 ( .A1(n5991), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n4890), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4882) );
  OAI211_X1 U6033 ( .C1(n5983), .C2(n5682), .A(n4883), .B(n4882), .ZN(n4885)
         );
  NOR2_X1 U6034 ( .A1(n5997), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4884)
         );
  AOI211_X1 U6035 ( .C1(n4887), .C2(n4886), .A(n4885), .B(n4884), .ZN(n4888)
         );
  OAI21_X1 U6036 ( .B1(n4902), .B2(n4889), .A(n4888), .ZN(U2826) );
  NOR2_X1 U6037 ( .A1(n4891), .A2(n4890), .ZN(n5990) );
  INV_X1 U6038 ( .A(REIP_REG_2__SCAN_IN), .ZN(n4898) );
  NAND2_X1 U6039 ( .A1(n4898), .A2(REIP_REG_1__SCAN_IN), .ZN(n4893) );
  NAND2_X1 U6040 ( .A1(n5991), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4892)
         );
  OAI21_X1 U6041 ( .B1(n5978), .B2(n4893), .A(n4892), .ZN(n4896) );
  NOR2_X1 U6042 ( .A1(n4894), .A2(n5996), .ZN(n4895) );
  AOI211_X1 U6043 ( .C1(n5993), .C2(EBX_REG_2__SCAN_IN), .A(n4896), .B(n4895), 
        .ZN(n4897) );
  OAI21_X1 U6044 ( .B1(n5990), .B2(n4898), .A(n4897), .ZN(n4900) );
  NOR2_X1 U6045 ( .A1(n5997), .A2(n6119), .ZN(n4899) );
  AOI211_X1 U6046 ( .C1(n5992), .C2(n6169), .A(n4900), .B(n4899), .ZN(n4901)
         );
  OAI21_X1 U6047 ( .B1(n4902), .B2(n6110), .A(n4901), .ZN(U2825) );
  NAND2_X1 U6048 ( .A1(n4926), .A2(n4903), .ZN(n4906) );
  NAND2_X1 U6049 ( .A1(n4904), .A2(n4927), .ZN(n4905) );
  XNOR2_X1 U6050 ( .A(n4906), .B(n4905), .ZN(n6131) );
  INV_X1 U6051 ( .A(n5912), .ZN(n6114) );
  NAND2_X1 U6052 ( .A1(n6131), .A2(n6114), .ZN(n4910) );
  INV_X1 U6053 ( .A(REIP_REG_9__SCAN_IN), .ZN(n4907) );
  NOR2_X1 U6054 ( .A1(n5585), .A2(n4907), .ZN(n6128) );
  NOR2_X1 U6055 ( .A1(n6118), .A2(n4919), .ZN(n4908) );
  AOI211_X1 U6056 ( .C1(n6109), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6128), 
        .B(n4908), .ZN(n4909) );
  OAI211_X1 U6057 ( .C1(n5591), .C2(n4911), .A(n4910), .B(n4909), .ZN(U2977)
         );
  INV_X1 U6058 ( .A(n4911), .ZN(n4912) );
  NAND2_X1 U6059 ( .A1(n4912), .A2(n5976), .ZN(n4918) );
  AOI22_X1 U6060 ( .A1(EBX_REG_9__SCAN_IN), .A2(n5993), .B1(
        REIP_REG_9__SCAN_IN), .B2(n5960), .ZN(n4913) );
  OAI211_X1 U6061 ( .C1(n5815), .C2(n3527), .A(n4913), .B(n5982), .ZN(n4916)
         );
  NOR2_X1 U6062 ( .A1(n5978), .A2(n4914), .ZN(n5962) );
  INV_X1 U6063 ( .A(n5962), .ZN(n4915) );
  NOR2_X1 U6064 ( .A1(n4915), .A2(REIP_REG_9__SCAN_IN), .ZN(n5961) );
  AOI211_X1 U6065 ( .C1(n6129), .C2(n5992), .A(n4916), .B(n5961), .ZN(n4917)
         );
  OAI211_X1 U6066 ( .C1(n4919), .C2(n5997), .A(n4918), .B(n4917), .ZN(U2818)
         );
  NAND2_X1 U6067 ( .A1(n4921), .A2(n4920), .ZN(n4922) );
  AND2_X1 U6068 ( .A1(n4983), .A2(n4922), .ZN(n5959) );
  INV_X1 U6069 ( .A(n5959), .ZN(n4953) );
  AOI22_X1 U6070 ( .A1(n5544), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n6014), .ZN(n4923) );
  OAI21_X1 U6071 ( .B1(n4953), .B2(n5862), .A(n4923), .ZN(U2881) );
  NAND2_X1 U6072 ( .A1(n5004), .A2(n4924), .ZN(n4930) );
  NAND2_X1 U6073 ( .A1(n4926), .A2(n4925), .ZN(n4928) );
  AND2_X1 U6074 ( .A1(n4928), .A2(n4927), .ZN(n4929) );
  XOR2_X1 U6075 ( .A(n4930), .B(n4929), .Z(n4958) );
  INV_X1 U6076 ( .A(n5687), .ZN(n5370) );
  OAI21_X1 U6077 ( .B1(n5370), .B2(n4934), .A(n6142), .ZN(n6130) );
  OAI21_X1 U6078 ( .B1(n4933), .B2(n4932), .A(n4986), .ZN(n5953) );
  INV_X1 U6079 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6442) );
  OAI22_X1 U6080 ( .A1(n5655), .A2(n5953), .B1(n6442), .B2(n5585), .ZN(n4936)
         );
  NAND2_X1 U6081 ( .A1(n4934), .A2(n6137), .ZN(n6134) );
  AOI221_X1 U6082 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n6515), .C2(n4799), .A(n6134), 
        .ZN(n4935) );
  AOI211_X1 U6083 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n6130), .A(n4936), .B(n4935), .ZN(n4937) );
  OAI21_X1 U6084 ( .B1(n4958), .B2(n5680), .A(n4937), .ZN(U3008) );
  INV_X1 U6085 ( .A(n4938), .ZN(n4939) );
  NAND2_X1 U6086 ( .A1(n4942), .A2(n4941), .ZN(n5031) );
  INV_X1 U6087 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4943) );
  NAND2_X1 U6088 ( .A1(n5581), .A2(n4943), .ZN(n4960) );
  NAND2_X1 U6089 ( .A1(n5230), .A2(n5028), .ZN(n5578) );
  XNOR2_X1 U6090 ( .A(n5581), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5120)
         );
  INV_X1 U6091 ( .A(n4944), .ZN(n4945) );
  NAND2_X1 U6092 ( .A1(n5875), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5034) );
  AND2_X1 U6093 ( .A1(n5037), .A2(n5034), .ZN(n5231) );
  NAND2_X1 U6094 ( .A1(n5578), .A2(n5231), .ZN(n4947) );
  XNOR2_X1 U6095 ( .A(n5581), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4946)
         );
  XNOR2_X1 U6096 ( .A(n4947), .B(n4946), .ZN(n5601) );
  NAND2_X1 U6097 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n4968), .ZN(n4972) );
  NOR2_X1 U6098 ( .A1(n4962), .A2(n4972), .ZN(n5048) );
  OAI21_X1 U6099 ( .B1(n5370), .B2(n5048), .A(n6127), .ZN(n5235) );
  NAND2_X1 U6100 ( .A1(n4948), .A2(n4974), .ZN(n4950) );
  INV_X1 U6101 ( .A(n5145), .ZN(n4949) );
  NAND2_X1 U6102 ( .A1(n4950), .A2(n4949), .ZN(n5465) );
  NAND2_X1 U6103 ( .A1(n6167), .A2(REIP_REG_15__SCAN_IN), .ZN(n5594) );
  OAI21_X1 U6104 ( .B1(n5655), .B2(n5465), .A(n5594), .ZN(n4951) );
  INV_X1 U6105 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6551) );
  INV_X1 U6106 ( .A(n5898), .ZN(n6122) );
  AND3_X1 U6107 ( .A1(n6551), .A2(n6122), .A3(n5048), .ZN(n5236) );
  AOI211_X1 U6108 ( .C1(n5235), .C2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n4951), .B(n5236), .ZN(n4952) );
  OAI21_X1 U6109 ( .B1(n5601), .B2(n5680), .A(n4952), .ZN(U3003) );
  OAI222_X1 U6110 ( .A1(n5953), .A2(n5535), .B1(n5532), .B2(n3036), .C1(n2945), 
        .C2(n4953), .ZN(U2849) );
  AOI22_X1 U6111 ( .A1(n6109), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6167), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n4954) );
  OAI21_X1 U6112 ( .B1(n6118), .B2(n4955), .A(n4954), .ZN(n4956) );
  AOI21_X1 U6113 ( .B1(n5959), .B2(n2946), .A(n4956), .ZN(n4957) );
  OAI21_X1 U6114 ( .B1(n4958), .B2(n5912), .A(n4957), .ZN(U2976) );
  NAND2_X1 U6115 ( .A1(n5230), .A2(n4959), .ZN(n5121) );
  NAND2_X1 U6116 ( .A1(n5121), .A2(n5120), .ZN(n4961) );
  NAND2_X1 U6117 ( .A1(n4961), .A2(n4960), .ZN(n4964) );
  XNOR2_X1 U6118 ( .A(n5581), .B(n4962), .ZN(n4963) );
  XNOR2_X1 U6119 ( .A(n4964), .B(n4963), .ZN(n5607) );
  NAND2_X1 U6120 ( .A1(n4965), .A2(n4972), .ZN(n4966) );
  OAI211_X1 U6121 ( .C1(n4967), .C2(n4968), .A(n6127), .B(n4966), .ZN(n5893)
         );
  NAND2_X1 U6122 ( .A1(n4943), .A2(n4968), .ZN(n5897) );
  INV_X1 U6123 ( .A(n5897), .ZN(n4970) );
  OAI221_X1 U6124 ( .B1(n5893), .B2(n4970), .C1(n5893), .C2(n4969), .A(
        INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4971) );
  INV_X1 U6125 ( .A(n4971), .ZN(n4980) );
  NOR3_X1 U6126 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5898), .A3(n4972), 
        .ZN(n4979) );
  INV_X1 U6127 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6448) );
  OR2_X1 U6128 ( .A1(n4973), .A2(n5139), .ZN(n4975) );
  NAND2_X1 U6129 ( .A1(n4975), .A2(n4974), .ZN(n5534) );
  INV_X1 U6130 ( .A(n5534), .ZN(n4976) );
  NAND2_X1 U6131 ( .A1(n6168), .A2(n4976), .ZN(n4977) );
  OAI21_X1 U6132 ( .B1(n6448), .B2(n5585), .A(n4977), .ZN(n4978) );
  NOR3_X1 U6133 ( .A1(n4980), .A2(n4979), .A3(n4978), .ZN(n4981) );
  OAI21_X1 U6134 ( .B1(n5607), .B2(n5680), .A(n4981), .ZN(U3004) );
  AND2_X1 U6135 ( .A1(n4983), .A2(n4982), .ZN(n4984) );
  OR2_X1 U6136 ( .A1(n4984), .A2(n5015), .ZN(n5012) );
  AOI21_X1 U6137 ( .B1(n4987), .B2(n4986), .A(n4985), .ZN(n6121) );
  AOI22_X1 U6138 ( .A1(n5511), .A2(n6121), .B1(n5509), .B2(EBX_REG_11__SCAN_IN), .ZN(n4988) );
  OAI21_X1 U6139 ( .B1(n5012), .B2(n2945), .A(n4988), .ZN(U2848) );
  AOI22_X1 U6140 ( .A1(n5544), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n6014), .ZN(n4989) );
  OAI21_X1 U6141 ( .B1(n5012), .B2(n5862), .A(n4989), .ZN(U2880) );
  INV_X1 U6142 ( .A(n5008), .ZN(n4998) );
  INV_X1 U6143 ( .A(n4990), .ZN(n4991) );
  NAND2_X1 U6144 ( .A1(n5962), .A2(n4991), .ZN(n5018) );
  OAI21_X1 U6145 ( .B1(n5978), .B2(n4993), .A(n4992), .ZN(n5938) );
  INV_X1 U6146 ( .A(n5938), .ZN(n4994) );
  AOI21_X1 U6147 ( .B1(n5017), .B2(n5018), .A(n4994), .ZN(n4997) );
  AOI22_X1 U6148 ( .A1(n5992), .A2(n6121), .B1(n5993), .B2(EBX_REG_11__SCAN_IN), .ZN(n4995) );
  OAI211_X1 U6149 ( .C1(n5815), .C2(n3559), .A(n4995), .B(n5982), .ZN(n4996)
         );
  AOI211_X1 U6150 ( .C1(n5958), .C2(n4998), .A(n4997), .B(n4996), .ZN(n4999)
         );
  OAI21_X1 U6151 ( .B1(n5820), .B2(n5012), .A(n4999), .ZN(U2816) );
  NAND2_X1 U6152 ( .A1(n5001), .A2(n5000), .ZN(n5003) );
  AND2_X1 U6153 ( .A1(n5003), .A2(n5002), .ZN(n5005) );
  NAND2_X1 U6154 ( .A1(n5005), .A2(n5004), .ZN(n5007) );
  XNOR2_X1 U6155 ( .A(n5581), .B(n6126), .ZN(n5006) );
  XNOR2_X1 U6156 ( .A(n5007), .B(n5006), .ZN(n6123) );
  NAND2_X1 U6157 ( .A1(n6123), .A2(n6114), .ZN(n5011) );
  NOR2_X1 U6158 ( .A1(n5585), .A2(n5017), .ZN(n6120) );
  NOR2_X1 U6159 ( .A1(n6118), .A2(n5008), .ZN(n5009) );
  AOI211_X1 U6160 ( .C1(n6109), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6120), 
        .B(n5009), .ZN(n5010) );
  OAI211_X1 U6161 ( .C1(n5591), .C2(n5012), .A(n5011), .B(n5010), .ZN(U2975)
         );
  OAI21_X1 U6162 ( .B1(n5015), .B2(n5014), .A(n5013), .ZN(n5130) );
  AOI22_X1 U6163 ( .A1(n5544), .A2(DATAI_12_), .B1(EAX_REG_12__SCAN_IN), .B2(
        n6014), .ZN(n5016) );
  OAI21_X1 U6164 ( .B1(n5130), .B2(n5862), .A(n5016), .ZN(U2879) );
  NOR2_X1 U6165 ( .A1(n5018), .A2(n5017), .ZN(n5939) );
  INV_X1 U6166 ( .A(n5939), .ZN(n5024) );
  NAND2_X1 U6167 ( .A1(n5991), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5019)
         );
  OAI211_X1 U6168 ( .C1(n5983), .C2(n5088), .A(n5982), .B(n5019), .ZN(n5022)
         );
  NOR2_X1 U6169 ( .A1(n5954), .A2(n5020), .ZN(n5021) );
  AOI211_X1 U6170 ( .C1(REIP_REG_12__SCAN_IN), .C2(n5938), .A(n5022), .B(n5021), .ZN(n5023) );
  OAI21_X1 U6171 ( .B1(n5024), .B2(REIP_REG_12__SCAN_IN), .A(n5023), .ZN(n5025) );
  AOI21_X1 U6172 ( .B1(n5958), .B2(n5133), .A(n5025), .ZN(n5026) );
  OAI21_X1 U6173 ( .B1(n5130), .B2(n5820), .A(n5026), .ZN(U2815) );
  NAND2_X1 U6174 ( .A1(n5581), .A2(n6551), .ZN(n5027) );
  INV_X1 U6175 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5579) );
  INV_X1 U6176 ( .A(n5251), .ZN(n5029) );
  NAND2_X1 U6177 ( .A1(n5031), .A2(n5030), .ZN(n5039) );
  OR2_X1 U6178 ( .A1(n5581), .A2(n6551), .ZN(n5232) );
  INV_X1 U6179 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5889) );
  INV_X1 U6180 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5678) );
  NAND3_X1 U6181 ( .A1(n5579), .A2(n5889), .A3(n5678), .ZN(n5032) );
  NAND2_X1 U6182 ( .A1(n5875), .A2(n5032), .ZN(n5033) );
  AND2_X1 U6183 ( .A1(n5232), .A2(n5033), .ZN(n5035) );
  AND2_X1 U6184 ( .A1(n5035), .A2(n5034), .ZN(n5036) );
  NAND2_X1 U6185 ( .A1(n5039), .A2(n5038), .ZN(n5041) );
  NAND2_X1 U6186 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5055) );
  NAND2_X1 U6187 ( .A1(n5581), .A2(n5055), .ZN(n5040) );
  NAND2_X2 U6188 ( .A1(n5041), .A2(n5040), .ZN(n5102) );
  NOR2_X1 U6189 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5658) );
  NOR2_X1 U6190 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5111) );
  INV_X1 U6191 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5342) );
  INV_X1 U6192 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5647) );
  NAND4_X1 U6193 ( .A1(n5658), .A2(n5111), .A3(n5342), .A4(n5647), .ZN(n5042)
         );
  NAND2_X1 U6194 ( .A1(n5875), .A2(n5042), .ZN(n5043) );
  NAND2_X1 U6195 ( .A1(n5102), .A2(n5043), .ZN(n5045) );
  AND2_X1 U6196 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5659) );
  AND2_X1 U6197 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5112) );
  AND2_X1 U6198 ( .A1(n5659), .A2(n5112), .ZN(n5254) );
  AND2_X1 U6199 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U6200 ( .A1(n5254), .A2(n5059), .ZN(n5095) );
  NAND2_X1 U6201 ( .A1(n5581), .A2(n5095), .ZN(n5044) );
  NAND2_X1 U6202 ( .A1(n5045), .A2(n5044), .ZN(n5047) );
  XNOR2_X1 U6203 ( .A(n5581), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5046)
         );
  OAI21_X1 U6204 ( .B1(n5047), .B2(n5046), .A(n5414), .ZN(n5289) );
  INV_X1 U6205 ( .A(n5289), .ZN(n5072) );
  NAND2_X1 U6206 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n5048), .ZN(n5240) );
  NOR2_X1 U6207 ( .A1(n5579), .A2(n5240), .ZN(n5051) );
  NAND2_X1 U6208 ( .A1(n5049), .A2(n5051), .ZN(n5062) );
  NAND2_X1 U6209 ( .A1(n5051), .A2(n5050), .ZN(n5064) );
  AOI22_X1 U6210 ( .A1(n5052), .A2(n5062), .B1(n6175), .B2(n5064), .ZN(n5053)
         );
  AND2_X1 U6211 ( .A1(n5054), .A2(n5053), .ZN(n5890) );
  INV_X1 U6212 ( .A(n5055), .ZN(n5066) );
  NAND2_X1 U6213 ( .A1(n5066), .A2(n5112), .ZN(n5339) );
  NAND2_X1 U6214 ( .A1(n5687), .A2(n5339), .ZN(n5056) );
  NAND2_X1 U6215 ( .A1(n5890), .A2(n5056), .ZN(n5668) );
  INV_X1 U6216 ( .A(n5659), .ZN(n5057) );
  AND2_X1 U6217 ( .A1(n5687), .A2(n5057), .ZN(n5058) );
  OR2_X1 U6218 ( .A1(n5668), .A2(n5058), .ZN(n5651) );
  INV_X1 U6219 ( .A(n6174), .ZN(n5060) );
  AOI21_X1 U6220 ( .B1(n5060), .B2(n5074), .A(n5059), .ZN(n5061) );
  NOR2_X1 U6221 ( .A1(n5651), .A2(n5061), .ZN(n5371) );
  INV_X1 U6222 ( .A(n5371), .ZN(n5099) );
  INV_X1 U6223 ( .A(n5062), .ZN(n5063) );
  NAND2_X1 U6224 ( .A1(n6174), .A2(n5063), .ZN(n5075) );
  OR2_X1 U6225 ( .A1(n5074), .A2(n5064), .ZN(n5065) );
  NAND2_X1 U6226 ( .A1(n5075), .A2(n5065), .ZN(n5885) );
  NAND2_X1 U6227 ( .A1(n5885), .A2(n5066), .ZN(n5113) );
  NOR2_X1 U6228 ( .A1(n5113), .A2(n5095), .ZN(n5364) );
  INV_X1 U6229 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5094) );
  AND2_X1 U6230 ( .A1(n5364), .A2(n5094), .ZN(n5098) );
  INV_X1 U6231 ( .A(n5497), .ZN(n5068) );
  AOI21_X1 U6232 ( .B1(n5068), .B2(n5270), .A(n5067), .ZN(n5069) );
  OR2_X1 U6233 ( .A1(n5069), .A2(n5092), .ZN(n5827) );
  NAND2_X1 U6234 ( .A1(n6167), .A2(REIP_REG_25__SCAN_IN), .ZN(n5286) );
  OAI21_X1 U6235 ( .B1(n5827), .B2(n5655), .A(n5286), .ZN(n5070) );
  AOI211_X1 U6236 ( .C1(n5099), .C2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5098), .B(n5070), .ZN(n5071) );
  OAI21_X1 U6237 ( .B1(n5072), .B2(n5680), .A(n5071), .ZN(U2993) );
  XNOR2_X2 U6238 ( .A(n5102), .B(n5073), .ZN(n5103) );
  XNOR2_X1 U6239 ( .A(n5103), .B(n5581), .ZN(n5576) );
  INV_X1 U6240 ( .A(n5890), .ZN(n5077) );
  AOI21_X1 U6241 ( .B1(n5075), .B2(n5074), .A(INSTADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n5076) );
  NOR2_X1 U6242 ( .A1(n5077), .A2(n5076), .ZN(n5679) );
  OAI21_X1 U6243 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5370), .A(n5679), 
        .ZN(n5115) );
  INV_X1 U6244 ( .A(n5105), .ZN(n5081) );
  NOR2_X1 U6245 ( .A1(n5079), .A2(n5078), .ZN(n5080) );
  AOI21_X1 U6246 ( .B1(n5081), .B2(n5078), .A(n5080), .ZN(n5454) );
  OR2_X1 U6247 ( .A1(n5528), .A2(n5454), .ZN(n5456) );
  INV_X1 U6248 ( .A(n5082), .ZN(n5083) );
  XNOR2_X1 U6249 ( .A(n5456), .B(n5083), .ZN(n5858) );
  INV_X1 U6250 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5084) );
  NOR2_X1 U6251 ( .A1(n5585), .A2(n5084), .ZN(n5572) );
  AOI21_X1 U6252 ( .B1(n6168), .B2(n5858), .A(n5572), .ZN(n5085) );
  OAI21_X1 U6253 ( .B1(n5113), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5085), 
        .ZN(n5086) );
  AOI21_X1 U6254 ( .B1(n5115), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5086), 
        .ZN(n5087) );
  OAI21_X1 U6255 ( .B1(n5576), .B2(n5680), .A(n5087), .ZN(U2999) );
  OAI222_X1 U6256 ( .A1(n5088), .A2(n5535), .B1(n5532), .B2(n5020), .C1(n2945), 
        .C2(n5130), .ZN(U2847) );
  AND2_X1 U6257 ( .A1(n5875), .A2(n6581), .ZN(n5547) );
  INV_X1 U6258 ( .A(n5547), .ZN(n5184) );
  NAND2_X1 U6259 ( .A1(n5581), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6260 ( .A1(n5184), .A2(n5183), .ZN(n5090) );
  NAND2_X1 U6261 ( .A1(n5581), .A2(n5094), .ZN(n5089) );
  XOR2_X1 U6262 ( .A(n5090), .B(n5549), .Z(n5320) );
  OR2_X1 U6263 ( .A1(n5092), .A2(n5091), .ZN(n5093) );
  AND2_X1 U6264 ( .A1(n5490), .A2(n5093), .ZN(n5322) );
  NAND2_X1 U6265 ( .A1(n6167), .A2(REIP_REG_26__SCAN_IN), .ZN(n5311) );
  INV_X1 U6266 ( .A(n5311), .ZN(n5097) );
  NOR4_X1 U6267 ( .A1(n5113), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n5095), 
        .A4(n5094), .ZN(n5096) );
  AOI211_X1 U6268 ( .C1(n6168), .C2(n5322), .A(n5097), .B(n5096), .ZN(n5101)
         );
  OAI21_X1 U6269 ( .B1(n5099), .B2(n5098), .A(INSTADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n5100) );
  OAI211_X1 U6270 ( .C1(n5320), .C2(n5680), .A(n5101), .B(n5100), .ZN(U2992)
         );
  OAI22_X1 U6271 ( .A1(n5103), .A2(n5581), .B1(n5102), .B2(n5073), .ZN(n5249)
         );
  XNOR2_X1 U6272 ( .A(n5581), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5248)
         );
  XNOR2_X1 U6273 ( .A(n5249), .B(n5248), .ZN(n5571) );
  NAND2_X1 U6274 ( .A1(n5106), .A2(n5432), .ZN(n5104) );
  OAI21_X1 U6275 ( .B1(n5106), .B2(n5105), .A(n5104), .ZN(n5109) );
  INV_X1 U6276 ( .A(n5107), .ZN(n5108) );
  XNOR2_X1 U6277 ( .A(n5109), .B(n5108), .ZN(n5510) );
  INV_X1 U6278 ( .A(REIP_REG_20__SCAN_IN), .ZN(n5110) );
  NOR2_X1 U6279 ( .A1(n5585), .A2(n5110), .ZN(n5566) );
  NOR3_X1 U6280 ( .A1(n5113), .A2(n5112), .A3(n5111), .ZN(n5114) );
  AOI211_X1 U6281 ( .C1(n6168), .C2(n5510), .A(n5566), .B(n5114), .ZN(n5117)
         );
  NAND2_X1 U6282 ( .A1(n5115), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5116) );
  OAI211_X1 U6283 ( .C1(n5571), .C2(n5680), .A(n5117), .B(n5116), .ZN(U2998)
         );
  OAI21_X1 U6284 ( .B1(n5119), .B2(n5118), .A(n5477), .ZN(n5136) );
  XNOR2_X1 U6285 ( .A(n5121), .B(n5120), .ZN(n5894) );
  NAND2_X1 U6286 ( .A1(n5894), .A2(n6114), .ZN(n5125) );
  INV_X1 U6287 ( .A(REIP_REG_13__SCAN_IN), .ZN(n5122) );
  NOR2_X1 U6288 ( .A1(n5585), .A2(n5122), .ZN(n5891) );
  NOR2_X1 U6289 ( .A1(n6118), .A2(n5947), .ZN(n5123) );
  AOI211_X1 U6290 ( .C1(n6109), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5891), 
        .B(n5123), .ZN(n5124) );
  OAI211_X1 U6291 ( .C1(n5591), .C2(n5136), .A(n5125), .B(n5124), .ZN(U2973)
         );
  INV_X1 U6292 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6022) );
  OAI222_X1 U6293 ( .A1(n5136), .A2(n5862), .B1(n5127), .B2(n5126), .C1(n6022), 
        .C2(n5421), .ZN(U2878) );
  INV_X1 U6294 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5129) );
  OAI21_X1 U6295 ( .B1(n5597), .B2(n5129), .A(n5128), .ZN(n5132) );
  NOR2_X1 U6296 ( .A1(n5130), .A2(n5591), .ZN(n5131) );
  AOI211_X1 U6297 ( .C1(n5593), .C2(n5133), .A(n5132), .B(n5131), .ZN(n5134)
         );
  OAI21_X1 U6298 ( .B1(n5135), .B2(n5912), .A(n5134), .ZN(U2974) );
  INV_X1 U6299 ( .A(n5136), .ZN(n5949) );
  NAND2_X1 U6300 ( .A1(n5138), .A2(n5137), .ZN(n5141) );
  INV_X1 U6301 ( .A(n5139), .ZN(n5140) );
  NAND2_X1 U6302 ( .A1(n5141), .A2(n5140), .ZN(n5945) );
  INV_X1 U6303 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5142) );
  OAI22_X1 U6304 ( .A1(n5535), .A2(n5945), .B1(n5142), .B2(n5532), .ZN(n5143)
         );
  AOI21_X1 U6305 ( .B1(n5949), .B2(n5537), .A(n5143), .ZN(n5144) );
  INV_X1 U6306 ( .A(n5144), .ZN(U2846) );
  OR2_X1 U6307 ( .A1(n5146), .A2(n5145), .ZN(n5147) );
  AND2_X1 U6308 ( .A1(n5526), .A2(n5147), .ZN(n5239) );
  INV_X1 U6309 ( .A(n5239), .ZN(n5151) );
  INV_X1 U6310 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6579) );
  INV_X1 U6311 ( .A(n5148), .ZN(n5150) );
  NAND2_X1 U6312 ( .A1(n5452), .A2(n5149), .ZN(n5522) );
  OAI21_X1 U6313 ( .B1(n5150), .B2(n5171), .A(n5522), .ZN(n5159) );
  OAI222_X1 U6314 ( .A1(n5151), .A2(n5535), .B1(n5532), .B2(n6579), .C1(n2945), 
        .C2(n5159), .ZN(U2843) );
  AOI21_X1 U6315 ( .B1(n5399), .B2(n5392), .A(n6488), .ZN(n5158) );
  NAND2_X1 U6316 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5398) );
  INV_X1 U6317 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5614) );
  AOI22_X1 U6318 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5614), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6583), .ZN(n5402) );
  NAND3_X1 U6319 ( .A1(n5399), .A2(n5152), .A3(n5157), .ZN(n5153) );
  OAI21_X1 U6320 ( .B1(n5398), .B2(n5402), .A(n5153), .ZN(n5154) );
  AOI21_X1 U6321 ( .B1(n5155), .B2(n5900), .A(n5154), .ZN(n5156) );
  OAI22_X1 U6322 ( .A1(n5158), .A2(n5157), .B1(n6488), .B2(n5156), .ZN(U3459)
         );
  INV_X1 U6323 ( .A(n5159), .ZN(n6013) );
  AND2_X1 U6324 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5160), .ZN(n5930) );
  INV_X1 U6325 ( .A(n5930), .ZN(n5164) );
  INV_X1 U6326 ( .A(n5459), .ZN(n5162) );
  NOR2_X1 U6327 ( .A1(n5162), .A2(n5161), .ZN(n5483) );
  NOR2_X1 U6328 ( .A1(n5978), .A2(REIP_REG_15__SCAN_IN), .ZN(n5466) );
  NOR2_X1 U6329 ( .A1(n5483), .A2(n5466), .ZN(n5163) );
  MUX2_X1 U6330 ( .A(n5164), .B(n5163), .S(REIP_REG_16__SCAN_IN), .Z(n5165) );
  OAI211_X1 U6331 ( .C1(n5815), .C2(n5166), .A(n5165), .B(n5982), .ZN(n5169)
         );
  AOI22_X1 U6332 ( .A1(n5992), .A2(n5239), .B1(n5993), .B2(EBX_REG_16__SCAN_IN), .ZN(n5167) );
  OAI21_X1 U6333 ( .B1(n5997), .B2(n5244), .A(n5167), .ZN(n5168) );
  AOI211_X1 U6334 ( .C1(n6013), .C2(n5976), .A(n5169), .B(n5168), .ZN(n5170)
         );
  INV_X1 U6335 ( .A(n5170), .ZN(U2811) );
  INV_X1 U6336 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5174) );
  AOI21_X1 U6337 ( .B1(n5173), .B2(n5172), .A(n5171), .ZN(n5599) );
  INV_X1 U6338 ( .A(n5599), .ZN(n5543) );
  OAI222_X1 U6339 ( .A1(n5465), .A2(n5535), .B1(n5174), .B2(n5532), .C1(n2945), 
        .C2(n5543), .ZN(U2844) );
  NAND2_X1 U6340 ( .A1(n5213), .A2(n5175), .ZN(n5177) );
  NAND2_X2 U6341 ( .A1(n5452), .A2(n5176), .ZN(n5500) );
  NOR2_X2 U6342 ( .A1(n5177), .A2(n5500), .ZN(n5282) );
  NAND2_X1 U6343 ( .A1(n5502), .A2(n5179), .ZN(n5427) );
  INV_X1 U6344 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6468) );
  NOR2_X1 U6345 ( .A1(n5585), .A2(n6468), .ZN(n5629) );
  NOR2_X1 U6346 ( .A1(n5597), .A2(n5181), .ZN(n5182) );
  AOI211_X1 U6347 ( .C1(n5199), .C2(n5593), .A(n5629), .B(n5182), .ZN(n5189)
         );
  INV_X1 U6348 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5640) );
  NOR2_X1 U6349 ( .A1(n5414), .A2(n5184), .ZN(n5294) );
  NAND2_X1 U6350 ( .A1(n5294), .A2(n5640), .ZN(n5185) );
  OAI21_X1 U6351 ( .B1(n5353), .B2(n5640), .A(n5185), .ZN(n5187) );
  XNOR2_X1 U6352 ( .A(n5187), .B(n5186), .ZN(n5635) );
  NAND2_X1 U6353 ( .A1(n5635), .A2(n6114), .ZN(n5188) );
  OAI211_X1 U6354 ( .C1(n5487), .C2(n5591), .A(n5189), .B(n5188), .ZN(U2958)
         );
  NOR3_X1 U6355 ( .A1(n6014), .A2(n5422), .A3(n5190), .ZN(n5191) );
  AOI22_X1 U6356 ( .A1(n6011), .A2(DATAI_12_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6014), .ZN(n5194) );
  NOR2_X2 U6357 ( .A1(n6014), .A2(n5192), .ZN(n6015) );
  NAND2_X1 U6358 ( .A1(n6015), .A2(DATAI_28_), .ZN(n5193) );
  OAI211_X1 U6359 ( .C1(n5487), .C2(n5862), .A(n5194), .B(n5193), .ZN(U2863)
         );
  NAND2_X1 U6360 ( .A1(n6468), .A2(REIP_REG_27__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U6361 ( .A1(n5492), .A2(n5195), .ZN(n5196) );
  NAND2_X1 U6362 ( .A1(n5430), .A2(n5196), .ZN(n5628) );
  AOI22_X1 U6363 ( .A1(n5993), .A2(EBX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n5991), .ZN(n5197) );
  OAI21_X1 U6364 ( .B1(n5628), .B2(n5983), .A(n5197), .ZN(n5198) );
  AOI21_X1 U6365 ( .B1(n5958), .B2(n5199), .A(n5198), .ZN(n5200) );
  OAI21_X1 U6366 ( .B1(n5814), .B2(n5201), .A(n5200), .ZN(n5202) );
  AOI21_X1 U6367 ( .B1(REIP_REG_28__SCAN_IN), .B2(n5439), .A(n5202), .ZN(n5203) );
  OAI21_X1 U6368 ( .B1(n5487), .B2(n5820), .A(n5203), .ZN(U2799) );
  INV_X1 U6369 ( .A(n5213), .ZN(n5204) );
  NOR2_X1 U6370 ( .A1(n5205), .A2(n5204), .ZN(n5313) );
  AND2_X1 U6371 ( .A1(n5313), .A2(n5502), .ZN(n5208) );
  INV_X1 U6372 ( .A(n5206), .ZN(n5207) );
  NOR2_X1 U6373 ( .A1(n5208), .A2(n5207), .ZN(n5209) );
  AOI22_X1 U6374 ( .A1(n6015), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6014), .ZN(n5212) );
  NAND2_X1 U6375 ( .A1(n6011), .A2(DATAI_11_), .ZN(n5211) );
  OAI211_X1 U6376 ( .C1(n5821), .C2(n5862), .A(n5212), .B(n5211), .ZN(U2864)
         );
  OR2_X1 U6377 ( .A1(n5502), .A2(n5213), .ZN(n5214) );
  AOI22_X1 U6378 ( .A1(n6011), .A2(DATAI_6_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n6014), .ZN(n5216) );
  NAND2_X1 U6379 ( .A1(n6015), .A2(DATAI_22_), .ZN(n5215) );
  OAI211_X1 U6380 ( .C1(n5304), .C2(n5862), .A(n5216), .B(n5215), .ZN(U2869)
         );
  INV_X1 U6381 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5222) );
  AND2_X1 U6382 ( .A1(n5506), .A2(n5217), .ZN(n5495) );
  INV_X1 U6383 ( .A(n5505), .ZN(n5220) );
  INV_X1 U6384 ( .A(n5218), .ZN(n5219) );
  AOI21_X1 U6385 ( .B1(n5506), .B2(n5220), .A(n5219), .ZN(n5221) );
  OR2_X1 U6386 ( .A1(n5495), .A2(n5221), .ZN(n5656) );
  OAI222_X1 U6387 ( .A1(n5222), .A2(n5532), .B1(n5535), .B2(n5656), .C1(n5304), 
        .C2(n2945), .ZN(U2837) );
  OAI22_X1 U6388 ( .A1(n5954), .A2(n5222), .B1(n5656), .B2(n5983), .ZN(n5224)
         );
  OAI22_X1 U6389 ( .A1(n5303), .A2(n5815), .B1(n5225), .B2(n5847), .ZN(n5223)
         );
  AOI211_X1 U6390 ( .C1(n5958), .C2(n5307), .A(n5224), .B(n5223), .ZN(n5228)
         );
  INV_X1 U6391 ( .A(n5836), .ZN(n5846) );
  AOI211_X1 U6392 ( .C1(n5225), .C2(n6457), .A(n5837), .B(n5846), .ZN(n5226)
         );
  INV_X1 U6393 ( .A(n5226), .ZN(n5227) );
  OAI211_X1 U6394 ( .C1(n5304), .C2(n5820), .A(n5228), .B(n5227), .ZN(U2805)
         );
  MUX2_X1 U6395 ( .A(n5579), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .S(n5581), 
        .Z(n5234) );
  NAND2_X1 U6396 ( .A1(n5230), .A2(n5229), .ZN(n5233) );
  XOR2_X1 U6397 ( .A(n5234), .B(n5252), .Z(n5247) );
  INV_X1 U6398 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6451) );
  OAI21_X1 U6399 ( .B1(n5236), .B2(n5235), .A(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n5237) );
  OAI21_X1 U6400 ( .B1(n5585), .B2(n6451), .A(n5237), .ZN(n5238) );
  AOI21_X1 U6401 ( .B1(n6168), .B2(n5239), .A(n5238), .ZN(n5242) );
  OR3_X1 U6402 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n5898), .A3(n5240), 
        .ZN(n5241) );
  OAI211_X1 U6403 ( .C1(n5247), .C2(n5680), .A(n5242), .B(n5241), .ZN(U3002)
         );
  AOI22_X1 U6404 ( .A1(n6109), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6167), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5243) );
  OAI21_X1 U6405 ( .B1(n6118), .B2(n5244), .A(n5243), .ZN(n5245) );
  AOI21_X1 U6406 ( .B1(n6013), .B2(n2946), .A(n5245), .ZN(n5246) );
  OAI21_X1 U6407 ( .B1(n5247), .B2(n5912), .A(n5246), .ZN(U2970) );
  AOI22_X1 U6408 ( .A1(n5249), .A2(n5248), .B1(n5875), .B2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5560) );
  XNOR2_X1 U6409 ( .A(n5581), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5559)
         );
  NAND2_X1 U6410 ( .A1(n5560), .A2(n5559), .ZN(n5558) );
  INV_X1 U6411 ( .A(n5558), .ZN(n5250) );
  NOR2_X1 U6412 ( .A1(n5581), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5301)
         );
  NAND2_X1 U6413 ( .A1(n5250), .A2(n5301), .ZN(n5335) );
  NAND2_X1 U6414 ( .A1(n5581), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5253) );
  NAND3_X1 U6415 ( .A1(n5881), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n5254), .ZN(n5255) );
  NAND2_X1 U6416 ( .A1(n5335), .A2(n5255), .ZN(n5256) );
  XNOR2_X1 U6417 ( .A(n5256), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5653)
         );
  NAND2_X1 U6418 ( .A1(n5264), .A2(n5257), .ZN(n5258) );
  INV_X1 U6419 ( .A(REIP_REG_23__SCAN_IN), .ZN(n5259) );
  OR2_X1 U6420 ( .A1(n5585), .A2(n5259), .ZN(n5648) );
  NAND2_X1 U6421 ( .A1(n6109), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5260)
         );
  OAI211_X1 U6422 ( .C1(n5844), .C2(n6118), .A(n5648), .B(n5260), .ZN(n5261)
         );
  AOI21_X1 U6423 ( .B1(n5863), .B2(n2946), .A(n5261), .ZN(n5262) );
  OAI21_X1 U6424 ( .B1(n5653), .B2(n5912), .A(n5262), .ZN(U2963) );
  OR2_X2 U6425 ( .A1(n5264), .A2(n5263), .ZN(n5284) );
  INV_X1 U6426 ( .A(n5284), .ZN(n5265) );
  AOI21_X1 U6427 ( .B1(n5267), .B2(n5266), .A(n5265), .ZN(n5350) );
  INV_X1 U6428 ( .A(n5350), .ZN(n5279) );
  AOI22_X1 U6429 ( .A1(n6011), .A2(DATAI_8_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6014), .ZN(n5269) );
  NAND2_X1 U6430 ( .A1(n6015), .A2(DATAI_24_), .ZN(n5268) );
  OAI211_X1 U6431 ( .C1(n5279), .C2(n5862), .A(n5269), .B(n5268), .ZN(U2867)
         );
  XNOR2_X1 U6432 ( .A(n5497), .B(n5270), .ZN(n5344) );
  AOI22_X1 U6433 ( .A1(n5344), .A2(n5511), .B1(EBX_REG_24__SCAN_IN), .B2(n5509), .ZN(n5271) );
  OAI21_X1 U6434 ( .B1(n5279), .B2(n2945), .A(n5271), .ZN(U2835) );
  INV_X1 U6435 ( .A(n5348), .ZN(n5277) );
  INV_X1 U6436 ( .A(n5344), .ZN(n5273) );
  NOR2_X1 U6437 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5325), .ZN(n5831) );
  AOI21_X1 U6438 ( .B1(n5993), .B2(EBX_REG_24__SCAN_IN), .A(n5831), .ZN(n5272)
         );
  OAI21_X1 U6439 ( .B1(n5273), .B2(n5983), .A(n5272), .ZN(n5276) );
  INV_X1 U6440 ( .A(REIP_REG_24__SCAN_IN), .ZN(n5326) );
  OAI22_X1 U6441 ( .A1(n5839), .A2(n5326), .B1(n5274), .B2(n5815), .ZN(n5275)
         );
  AOI211_X1 U6442 ( .C1(n5958), .C2(n5277), .A(n5276), .B(n5275), .ZN(n5278)
         );
  OAI21_X1 U6443 ( .B1(n5279), .B2(n5820), .A(n5278), .ZN(U2803) );
  INV_X1 U6444 ( .A(n5280), .ZN(n5281) );
  INV_X1 U6445 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5287) );
  OAI21_X1 U6446 ( .B1(n5597), .B2(n5287), .A(n5286), .ZN(n5288) );
  AOI21_X1 U6447 ( .B1(n5826), .B2(n5593), .A(n5288), .ZN(n5291) );
  NAND2_X1 U6448 ( .A1(n5289), .A2(n6114), .ZN(n5290) );
  OAI211_X1 U6449 ( .C1(n5310), .C2(n5591), .A(n5291), .B(n5290), .ZN(U2961)
         );
  AOI22_X1 U6450 ( .A1(n6015), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6014), .ZN(n5293) );
  NAND2_X1 U6451 ( .A1(n6011), .A2(DATAI_9_), .ZN(n5292) );
  OAI211_X1 U6452 ( .C1(n5310), .C2(n5862), .A(n5293), .B(n5292), .ZN(U2866)
         );
  INV_X1 U6453 ( .A(n5353), .ZN(n5295) );
  NOR2_X1 U6454 ( .A1(n5295), .A2(n5294), .ZN(n5296) );
  XNOR2_X1 U6455 ( .A(n5296), .B(n5640), .ZN(n5646) );
  INV_X1 U6456 ( .A(n5821), .ZN(n5299) );
  INV_X1 U6457 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6464) );
  NOR2_X1 U6458 ( .A1(n5585), .A2(n6464), .ZN(n5638) );
  AOI21_X1 U6459 ( .B1(n6109), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5638), 
        .ZN(n5297) );
  OAI21_X1 U6460 ( .B1(n5813), .B2(n6118), .A(n5297), .ZN(n5298) );
  AOI21_X1 U6461 ( .B1(n5299), .B2(n2946), .A(n5298), .ZN(n5300) );
  OAI21_X1 U6462 ( .B1(n5646), .B2(n5912), .A(n5300), .ZN(U2959) );
  OAI21_X1 U6463 ( .B1(n5875), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5558), 
        .ZN(n5337) );
  AOI21_X1 U6464 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5581), .A(n5301), 
        .ZN(n5302) );
  XNOR2_X1 U6465 ( .A(n5337), .B(n5302), .ZN(n5663) );
  OR2_X1 U6466 ( .A1(n5585), .A2(n5225), .ZN(n5654) );
  OAI21_X1 U6467 ( .B1(n5597), .B2(n5303), .A(n5654), .ZN(n5306) );
  NOR2_X1 U6468 ( .A1(n5304), .A2(n5591), .ZN(n5305) );
  AOI211_X1 U6469 ( .C1(n5593), .C2(n5307), .A(n5306), .B(n5305), .ZN(n5308)
         );
  OAI21_X1 U6470 ( .B1(n5663), .B2(n5912), .A(n5308), .ZN(U2964) );
  OAI222_X1 U6471 ( .A1(n5310), .A2(n2945), .B1(n5532), .B2(n5309), .C1(n5827), 
        .C2(n5535), .ZN(U2834) );
  OAI21_X1 U6472 ( .B1(n5597), .B2(n5312), .A(n5311), .ZN(n5318) );
  NAND2_X1 U6473 ( .A1(n5502), .A2(n5313), .ZN(n5314) );
  OAI21_X2 U6474 ( .B1(n5316), .B2(n5315), .A(n5314), .ZN(n5334) );
  NOR2_X1 U6475 ( .A1(n5334), .A2(n5591), .ZN(n5317) );
  AOI211_X1 U6476 ( .C1(n5330), .C2(n5593), .A(n5318), .B(n5317), .ZN(n5319)
         );
  OAI21_X1 U6477 ( .B1(n5320), .B2(n5912), .A(n5319), .ZN(U2960) );
  AOI22_X1 U6478 ( .A1(n5322), .A2(n5511), .B1(n5509), .B2(EBX_REG_26__SCAN_IN), .ZN(n5321) );
  OAI21_X1 U6479 ( .B1(n5334), .B2(n2945), .A(n5321), .ZN(U2833) );
  INV_X1 U6480 ( .A(n5322), .ZN(n5324) );
  AOI22_X1 U6481 ( .A1(EBX_REG_26__SCAN_IN), .A2(n5993), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n5991), .ZN(n5323) );
  OAI21_X1 U6482 ( .B1(n5983), .B2(n5324), .A(n5323), .ZN(n5329) );
  NOR2_X1 U6483 ( .A1(n5326), .A2(n5325), .ZN(n5825) );
  AOI21_X1 U6484 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5825), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5327) );
  NOR2_X1 U6485 ( .A1(n5327), .A2(n5816), .ZN(n5328) );
  AOI211_X1 U6486 ( .C1(n5958), .C2(n5330), .A(n5329), .B(n5328), .ZN(n5331)
         );
  OAI21_X1 U6487 ( .B1(n5334), .B2(n5820), .A(n5331), .ZN(U2801) );
  AOI22_X1 U6488 ( .A1(n6011), .A2(DATAI_10_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6014), .ZN(n5333) );
  NAND2_X1 U6489 ( .A1(n6015), .A2(DATAI_26_), .ZN(n5332) );
  OAI211_X1 U6490 ( .C1(n5334), .C2(n5862), .A(n5333), .B(n5332), .ZN(U2865)
         );
  NAND3_X1 U6491 ( .A1(n5581), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5336) );
  XNOR2_X1 U6492 ( .A(n5338), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5352)
         );
  NOR2_X1 U6493 ( .A1(n5585), .A2(n5326), .ZN(n5346) );
  INV_X1 U6494 ( .A(n5339), .ZN(n5340) );
  AND2_X1 U6495 ( .A1(n5885), .A2(n5340), .ZN(n5657) );
  NAND3_X1 U6496 ( .A1(n5657), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n5659), .ZN(n5341) );
  AOI21_X1 U6497 ( .B1(n5342), .B2(n5341), .A(n5371), .ZN(n5343) );
  AOI211_X1 U6498 ( .C1(n6168), .C2(n5344), .A(n5346), .B(n5343), .ZN(n5345)
         );
  OAI21_X1 U6499 ( .B1(n5352), .B2(n5680), .A(n5345), .ZN(U2994) );
  AOI21_X1 U6500 ( .B1(n6109), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5346), 
        .ZN(n5347) );
  OAI21_X1 U6501 ( .B1(n5348), .B2(n6118), .A(n5347), .ZN(n5349) );
  AOI21_X1 U6502 ( .B1(n5350), .B2(n2946), .A(n5349), .ZN(n5351) );
  OAI21_X1 U6503 ( .B1(n5352), .B2(n5912), .A(n5351), .ZN(U2962) );
  NAND2_X1 U6504 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5369) );
  NOR2_X2 U6505 ( .A1(n5353), .A2(n5369), .ZN(n5551) );
  NOR2_X1 U6506 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5548) );
  INV_X1 U6507 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6552) );
  NAND3_X1 U6508 ( .A1(n5547), .A2(n5548), .A3(n6552), .ZN(n5413) );
  INV_X1 U6509 ( .A(n5413), .ZN(n5354) );
  OAI22_X1 U6510 ( .A1(n5551), .A2(n5354), .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5549), .ZN(n5355) );
  XOR2_X1 U6511 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .B(n5355), .Z(n5382) );
  INV_X1 U6512 ( .A(n5430), .ZN(n5358) );
  INV_X1 U6513 ( .A(n5359), .ZN(n5356) );
  OAI211_X1 U6514 ( .C1(n5358), .C2(n5078), .A(n5357), .B(n5356), .ZN(n5363)
         );
  OAI211_X1 U6515 ( .C1(n5361), .C2(n5430), .A(n5360), .B(n5359), .ZN(n5362)
         );
  NAND2_X1 U6516 ( .A1(n5363), .A2(n5362), .ZN(n5409) );
  INV_X1 U6517 ( .A(n5409), .ZN(n5367) );
  NAND2_X1 U6518 ( .A1(n6167), .A2(REIP_REG_30__SCAN_IN), .ZN(n5377) );
  INV_X1 U6519 ( .A(n5377), .ZN(n5366) );
  AND2_X1 U6520 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5368) );
  NAND2_X1 U6521 ( .A1(n5364), .A2(n5368), .ZN(n5637) );
  NOR2_X1 U6522 ( .A1(n5637), .A2(n5369), .ZN(n5611) );
  INV_X1 U6523 ( .A(n5611), .ZN(n5623) );
  NOR3_X1 U6524 ( .A1(n5623), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n6552), 
        .ZN(n5365) );
  AOI211_X1 U6525 ( .C1(n5367), .C2(n6168), .A(n5366), .B(n5365), .ZN(n5374)
         );
  NAND2_X1 U6526 ( .A1(n5371), .A2(n5368), .ZN(n5642) );
  OR2_X1 U6527 ( .A1(n5642), .A2(n5369), .ZN(n5372) );
  NAND2_X1 U6528 ( .A1(n5371), .A2(n5370), .ZN(n5643) );
  AND2_X1 U6529 ( .A1(n5372), .A2(n5643), .ZN(n5625) );
  OAI211_X1 U6530 ( .C1(n5625), .C2(n6552), .A(INSTADDRPOINTER_REG_30__SCAN_IN), .B(n5643), .ZN(n5373) );
  OAI211_X1 U6531 ( .C1(n5382), .C2(n5680), .A(n5374), .B(n5373), .ZN(U2988)
         );
  XOR2_X1 U6532 ( .A(n5426), .B(n5376), .Z(n5406) );
  NAND2_X1 U6533 ( .A1(n5387), .A2(n5593), .ZN(n5378) );
  OAI211_X1 U6534 ( .C1(n5597), .C2(n5379), .A(n5378), .B(n5377), .ZN(n5380)
         );
  AOI21_X1 U6535 ( .B1(n5406), .B2(n2946), .A(n5380), .ZN(n5381) );
  OAI21_X1 U6536 ( .B1(n5912), .B2(n5382), .A(n5381), .ZN(U2956) );
  NAND2_X1 U6537 ( .A1(n5406), .A2(n5976), .ZN(n5389) );
  AOI22_X1 U6538 ( .A1(n5993), .A2(EBX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n5991), .ZN(n5383) );
  OAI21_X1 U6539 ( .B1(n5409), .B2(n5983), .A(n5383), .ZN(n5386) );
  NOR3_X1 U6540 ( .A1(n5384), .A2(REIP_REG_30__SCAN_IN), .A3(n6470), .ZN(n5385) );
  AOI211_X1 U6541 ( .C1(n5387), .C2(n5958), .A(n5386), .B(n5385), .ZN(n5388)
         );
  OAI211_X1 U6542 ( .C1(n5390), .C2(n6473), .A(n5389), .B(n5388), .ZN(U2797)
         );
  INV_X1 U6543 ( .A(n5391), .ZN(n5393) );
  NAND3_X1 U6544 ( .A1(n5394), .A2(n5393), .A3(n5392), .ZN(n5395) );
  OAI211_X1 U6545 ( .C1(n5693), .C2(n5397), .A(n5396), .B(n5395), .ZN(n6370)
         );
  INV_X1 U6546 ( .A(n5398), .ZN(n5401) );
  AOI222_X1 U6547 ( .A1(n6370), .A2(n5900), .B1(n5402), .B2(n5401), .C1(n5400), 
        .C2(n5399), .ZN(n5405) );
  OAI22_X1 U6548 ( .A1(n6488), .A2(n5405), .B1(n5404), .B2(n5403), .ZN(U3460)
         );
  INV_X1 U6549 ( .A(n5406), .ZN(n5411) );
  AOI22_X1 U6550 ( .A1(n6011), .A2(DATAI_14_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6014), .ZN(n5408) );
  NAND2_X1 U6551 ( .A1(n6015), .A2(DATAI_30_), .ZN(n5407) );
  OAI211_X1 U6552 ( .C1(n5411), .C2(n5862), .A(n5408), .B(n5407), .ZN(U2861)
         );
  INV_X1 U6553 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5410) );
  OAI222_X1 U6554 ( .A1(n2945), .A2(n5411), .B1(n5532), .B2(n5410), .C1(n5409), 
        .C2(n5535), .ZN(U2829) );
  OAI22_X1 U6555 ( .A1(n5608), .A2(n5535), .B1(n5412), .B2(n5532), .ZN(U2828)
         );
  AND2_X1 U6556 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5610) );
  NOR3_X1 U6557 ( .A1(n5414), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5413), 
        .ZN(n5415) );
  AOI21_X1 U6558 ( .B1(n5551), .B2(n5610), .A(n5415), .ZN(n5416) );
  XNOR2_X1 U6559 ( .A(n5416), .B(n5614), .ZN(n5619) );
  NAND2_X1 U6560 ( .A1(n6167), .A2(REIP_REG_31__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U6561 ( .A1(n6109), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5417)
         );
  OAI211_X1 U6562 ( .C1(n5418), .C2(n6118), .A(n5613), .B(n5417), .ZN(n5419)
         );
  AOI21_X1 U6563 ( .B1(n5423), .B2(n2946), .A(n5419), .ZN(n5420) );
  OAI21_X1 U6564 ( .B1(n5619), .B2(n5912), .A(n5420), .ZN(U2955) );
  NAND3_X1 U6565 ( .A1(n5423), .A2(n5422), .A3(n5421), .ZN(n5425) );
  AOI22_X1 U6566 ( .A1(n6015), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6014), .ZN(n5424) );
  NAND2_X1 U6567 ( .A1(n5425), .A2(n5424), .ZN(U2860) );
  AOI21_X1 U6568 ( .B1(n5428), .B2(n5427), .A(n5426), .ZN(n5556) );
  INV_X1 U6569 ( .A(n5556), .ZN(n5541) );
  AOI22_X1 U6570 ( .A1(n5993), .A2(EBX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n5991), .ZN(n5436) );
  OAI211_X1 U6571 ( .C1(n5432), .C2(n5431), .A(n5430), .B(n5429), .ZN(n5433)
         );
  AND2_X1 U6572 ( .A1(n5434), .A2(n5433), .ZN(n5621) );
  NAND2_X1 U6573 ( .A1(n5621), .A2(n5992), .ZN(n5435) );
  OAI211_X1 U6574 ( .C1(n5997), .C2(n5554), .A(n5436), .B(n5435), .ZN(n5438)
         );
  AOI211_X1 U6575 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5439), .A(n5438), .B(n5437), .ZN(n5440) );
  OAI21_X1 U6576 ( .B1(n5541), .B2(n5820), .A(n5440), .ZN(U2798) );
  XOR2_X1 U6577 ( .A(n5441), .B(n5500), .Z(n5869) );
  INV_X1 U6578 ( .A(n5869), .ZN(n5513) );
  INV_X1 U6579 ( .A(n5510), .ZN(n5442) );
  OAI22_X1 U6580 ( .A1(n5954), .A2(n5443), .B1(n5442), .B2(n5983), .ZN(n5448)
         );
  INV_X1 U6581 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6453) );
  NOR2_X1 U6582 ( .A1(n5084), .A2(n6453), .ZN(n5854) );
  INV_X1 U6583 ( .A(n5853), .ZN(n5444) );
  AOI21_X1 U6584 ( .B1(n5854), .B2(n5444), .A(REIP_REG_20__SCAN_IN), .ZN(n5446) );
  OAI22_X1 U6585 ( .A1(n5446), .A2(n5847), .B1(n5445), .B2(n5815), .ZN(n5447)
         );
  AOI211_X1 U6586 ( .C1(n5958), .C2(n5565), .A(n5448), .B(n5447), .ZN(n5449)
         );
  OAI21_X1 U6587 ( .B1(n5513), .B2(n5820), .A(n5449), .ZN(U2807) );
  AND2_X1 U6588 ( .A1(n5452), .A2(n5450), .ZN(n5524) );
  NAND2_X1 U6589 ( .A1(n5452), .A2(n5451), .ZN(n5515) );
  OAI21_X1 U6590 ( .B1(n5524), .B2(n5453), .A(n5515), .ZN(n6004) );
  NAND2_X1 U6591 ( .A1(n5528), .A2(n5454), .ZN(n5455) );
  AND2_X1 U6592 ( .A1(n5456), .A2(n5455), .ZN(n5675) );
  INV_X1 U6593 ( .A(n5675), .ZN(n5520) );
  OAI22_X1 U6594 ( .A1(n5954), .A2(n5457), .B1(n5983), .B2(n5520), .ZN(n5462)
         );
  NAND2_X1 U6595 ( .A1(n5459), .A2(n5458), .ZN(n5931) );
  AOI21_X1 U6596 ( .B1(n5991), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5956), 
        .ZN(n5460) );
  OAI221_X1 U6597 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5853), .C1(n6453), .C2(
        n5931), .A(n5460), .ZN(n5461) );
  AOI211_X1 U6598 ( .C1(n5958), .C2(n5586), .A(n5462), .B(n5461), .ZN(n5463)
         );
  OAI21_X1 U6599 ( .B1(n6004), .B2(n5820), .A(n5463), .ZN(U2809) );
  AOI21_X1 U6600 ( .B1(n5991), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5956), 
        .ZN(n5464) );
  OAI21_X1 U6601 ( .B1(n5983), .B2(n5465), .A(n5464), .ZN(n5471) );
  INV_X1 U6602 ( .A(n5466), .ZN(n5468) );
  AOI22_X1 U6603 ( .A1(EBX_REG_15__SCAN_IN), .A2(n5993), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5483), .ZN(n5467) );
  OAI21_X1 U6604 ( .B1(n5469), .B2(n5468), .A(n5467), .ZN(n5470) );
  AOI211_X1 U6605 ( .C1(n5592), .C2(n5958), .A(n5471), .B(n5470), .ZN(n5472)
         );
  OAI21_X1 U6606 ( .B1(n5543), .B2(n5820), .A(n5472), .ZN(U2812) );
  INV_X1 U6607 ( .A(n5473), .ZN(n5475) );
  NOR2_X1 U6608 ( .A1(n5475), .A2(n5474), .ZN(n5478) );
  AOI21_X1 U6609 ( .B1(n5478), .B2(n5477), .A(n5476), .ZN(n5605) );
  INV_X1 U6610 ( .A(n5605), .ZN(n5546) );
  NAND2_X1 U6611 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5939), .ZN(n5941) );
  OAI21_X1 U6612 ( .B1(n5122), .B2(n5941), .A(n6448), .ZN(n5484) );
  NAND2_X1 U6613 ( .A1(n5991), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5479)
         );
  OAI211_X1 U6614 ( .C1(n5983), .C2(n5534), .A(n5982), .B(n5479), .ZN(n5480)
         );
  AOI21_X1 U6615 ( .B1(n5993), .B2(EBX_REG_14__SCAN_IN), .A(n5480), .ZN(n5481)
         );
  OAI21_X1 U6616 ( .B1(n5997), .B2(n5603), .A(n5481), .ZN(n5482) );
  AOI21_X1 U6617 ( .B1(n5484), .B2(n5483), .A(n5482), .ZN(n5485) );
  OAI21_X1 U6618 ( .B1(n5546), .B2(n5820), .A(n5485), .ZN(U2813) );
  AOI22_X1 U6619 ( .A1(n5621), .A2(n5511), .B1(n5509), .B2(EBX_REG_29__SCAN_IN), .ZN(n5486) );
  OAI21_X1 U6620 ( .B1(n5541), .B2(n2945), .A(n5486), .ZN(U2830) );
  OAI222_X1 U6621 ( .A1(n5488), .A2(n5532), .B1(n5535), .B2(n5628), .C1(n5487), 
        .C2(n2945), .ZN(U2831) );
  INV_X1 U6622 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U6623 ( .A1(n5490), .A2(n5489), .ZN(n5491) );
  NAND2_X1 U6624 ( .A1(n5492), .A2(n5491), .ZN(n5819) );
  OAI222_X1 U6625 ( .A1(n2945), .A2(n5821), .B1(n5532), .B2(n5493), .C1(n5819), 
        .C2(n5535), .ZN(U2832) );
  INV_X1 U6626 ( .A(n5863), .ZN(n5499) );
  INV_X1 U6627 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5498) );
  OR2_X1 U6628 ( .A1(n5495), .A2(n5494), .ZN(n5496) );
  NAND2_X1 U6629 ( .A1(n5497), .A2(n5496), .ZN(n5838) );
  OAI222_X1 U6630 ( .A1(n2945), .A2(n5499), .B1(n5532), .B2(n5498), .C1(n5838), 
        .C2(n5535), .ZN(U2836) );
  INV_X1 U6631 ( .A(n5500), .ZN(n5514) );
  NAND2_X1 U6632 ( .A1(n5514), .A2(n5501), .ZN(n5503) );
  AOI21_X1 U6633 ( .B1(n5504), .B2(n5503), .A(n5502), .ZN(n5866) );
  INV_X1 U6634 ( .A(n5866), .ZN(n5508) );
  XNOR2_X1 U6635 ( .A(n5506), .B(n5505), .ZN(n5849) );
  INV_X1 U6636 ( .A(n5849), .ZN(n5507) );
  OAI222_X1 U6637 ( .A1(n5508), .A2(n2945), .B1(n5535), .B2(n5507), .C1(n5532), 
        .C2(n3076), .ZN(U2838) );
  AOI22_X1 U6638 ( .A1(n5511), .A2(n5510), .B1(EBX_REG_20__SCAN_IN), .B2(n5509), .ZN(n5512) );
  OAI21_X1 U6639 ( .B1(n5513), .B2(n2945), .A(n5512), .ZN(U2839) );
  AOI21_X1 U6640 ( .B1(n5516), .B2(n5515), .A(n5514), .ZN(n5872) );
  INV_X1 U6641 ( .A(n5872), .ZN(n5519) );
  INV_X1 U6642 ( .A(n5858), .ZN(n5518) );
  OAI222_X1 U6643 ( .A1(n5519), .A2(n2945), .B1(n5535), .B2(n5518), .C1(n5517), 
        .C2(n5532), .ZN(U2840) );
  OAI222_X1 U6644 ( .A1(n5520), .A2(n5535), .B1(n5532), .B2(n5457), .C1(n2945), 
        .C2(n6004), .ZN(U2841) );
  AND2_X1 U6645 ( .A1(n5522), .A2(n5521), .ZN(n5523) );
  NAND2_X1 U6646 ( .A1(n5526), .A2(n5525), .ZN(n5527) );
  AND2_X1 U6647 ( .A1(n5528), .A2(n5527), .ZN(n5934) );
  INV_X1 U6648 ( .A(n5934), .ZN(n5529) );
  INV_X1 U6649 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6623) );
  OAI22_X1 U6650 ( .A1(n5535), .A2(n5529), .B1(n6623), .B2(n5532), .ZN(n5530)
         );
  AOI21_X1 U6651 ( .B1(n6008), .B2(n5537), .A(n5530), .ZN(n5531) );
  INV_X1 U6652 ( .A(n5531), .ZN(U2842) );
  OAI22_X1 U6653 ( .A1(n5535), .A2(n5534), .B1(n5533), .B2(n5532), .ZN(n5536)
         );
  AOI21_X1 U6654 ( .B1(n5605), .B2(n5537), .A(n5536), .ZN(n5538) );
  INV_X1 U6655 ( .A(n5538), .ZN(U2845) );
  AOI22_X1 U6656 ( .A1(n6011), .A2(DATAI_13_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6014), .ZN(n5540) );
  NAND2_X1 U6657 ( .A1(n6015), .A2(DATAI_29_), .ZN(n5539) );
  OAI211_X1 U6658 ( .C1(n5541), .C2(n5862), .A(n5540), .B(n5539), .ZN(U2862)
         );
  AOI22_X1 U6659 ( .A1(n5544), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6014), .ZN(n5542) );
  OAI21_X1 U6660 ( .B1(n5543), .B2(n5862), .A(n5542), .ZN(U2876) );
  AOI22_X1 U6661 ( .A1(n5544), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n6014), .ZN(n5545) );
  OAI21_X1 U6662 ( .B1(n5546), .B2(n5862), .A(n5545), .ZN(U2877) );
  AND3_X1 U6663 ( .A1(n5549), .A2(n5548), .A3(n5547), .ZN(n5550) );
  OR2_X1 U6664 ( .A1(n5551), .A2(n5550), .ZN(n5552) );
  XNOR2_X1 U6665 ( .A(n5552), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5627)
         );
  NOR2_X1 U6666 ( .A1(n5585), .A2(n6470), .ZN(n5620) );
  AOI21_X1 U6667 ( .B1(n6109), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5620), 
        .ZN(n5553) );
  OAI21_X1 U6668 ( .B1(n5554), .B2(n6118), .A(n5553), .ZN(n5555) );
  AOI21_X1 U6669 ( .B1(n5556), .B2(n2946), .A(n5555), .ZN(n5557) );
  OAI21_X1 U6670 ( .B1(n5627), .B2(n5912), .A(n5557), .ZN(U2957) );
  OAI21_X1 U6671 ( .B1(n5560), .B2(n5559), .A(n5558), .ZN(n5561) );
  INV_X1 U6672 ( .A(n5561), .ZN(n5670) );
  NAND2_X1 U6673 ( .A1(n6167), .A2(REIP_REG_21__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U6674 ( .A1(n6109), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5562)
         );
  OAI211_X1 U6675 ( .C1(n5852), .C2(n6118), .A(n5664), .B(n5562), .ZN(n5563)
         );
  AOI21_X1 U6676 ( .B1(n5866), .B2(n2946), .A(n5563), .ZN(n5564) );
  OAI21_X1 U6677 ( .B1(n5670), .B2(n5912), .A(n5564), .ZN(U2965) );
  INV_X1 U6678 ( .A(n5565), .ZN(n5568) );
  AOI21_X1 U6679 ( .B1(n6109), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5566), 
        .ZN(n5567) );
  OAI21_X1 U6680 ( .B1(n6118), .B2(n5568), .A(n5567), .ZN(n5569) );
  AOI21_X1 U6681 ( .B1(n5869), .B2(n2946), .A(n5569), .ZN(n5570) );
  OAI21_X1 U6682 ( .B1(n5571), .B2(n5912), .A(n5570), .ZN(U2966) );
  AOI21_X1 U6683 ( .B1(n6109), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5572), 
        .ZN(n5573) );
  OAI21_X1 U6684 ( .B1(n5861), .B2(n6118), .A(n5573), .ZN(n5574) );
  AOI21_X1 U6685 ( .B1(n5872), .B2(n2946), .A(n5574), .ZN(n5575) );
  OAI21_X1 U6686 ( .B1(n5576), .B2(n5912), .A(n5575), .ZN(U2967) );
  NAND2_X1 U6687 ( .A1(n5578), .A2(n5577), .ZN(n5583) );
  NAND2_X1 U6688 ( .A1(n5579), .A2(n5889), .ZN(n5580) );
  OR2_X1 U6689 ( .A1(n5581), .A2(n5580), .ZN(n5582) );
  NOR2_X1 U6690 ( .A1(n5583), .A2(n5582), .ZN(n5879) );
  NOR2_X1 U6691 ( .A1(n5881), .A2(n5879), .ZN(n5584) );
  XNOR2_X1 U6692 ( .A(n5584), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5671)
         );
  NAND2_X1 U6693 ( .A1(n5671), .A2(n6114), .ZN(n5590) );
  NOR2_X1 U6694 ( .A1(n5585), .A2(n6453), .ZN(n5674) );
  INV_X1 U6695 ( .A(n5586), .ZN(n5587) );
  NOR2_X1 U6696 ( .A1(n5587), .A2(n6118), .ZN(n5588) );
  AOI211_X1 U6697 ( .C1(n6109), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5674), 
        .B(n5588), .ZN(n5589) );
  OAI211_X1 U6698 ( .C1(n5591), .C2(n6004), .A(n5590), .B(n5589), .ZN(U2968)
         );
  INV_X1 U6699 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U6700 ( .A1(n5593), .A2(n5592), .ZN(n5595) );
  OAI211_X1 U6701 ( .C1(n5597), .C2(n5596), .A(n5595), .B(n5594), .ZN(n5598)
         );
  AOI21_X1 U6702 ( .B1(n5599), .B2(n2946), .A(n5598), .ZN(n5600) );
  OAI21_X1 U6703 ( .B1(n5601), .B2(n5912), .A(n5600), .ZN(U2971) );
  AOI22_X1 U6704 ( .A1(n6109), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6167), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5602) );
  OAI21_X1 U6705 ( .B1(n6118), .B2(n5603), .A(n5602), .ZN(n5604) );
  AOI21_X1 U6706 ( .B1(n5605), .B2(n2946), .A(n5604), .ZN(n5606) );
  OAI21_X1 U6707 ( .B1(n5607), .B2(n5912), .A(n5606), .ZN(U2972) );
  INV_X1 U6708 ( .A(n5608), .ZN(n5617) );
  INV_X1 U6709 ( .A(n5610), .ZN(n5609) );
  AOI21_X1 U6710 ( .B1(n5687), .B2(n5609), .A(n5625), .ZN(n5615) );
  NAND3_X1 U6711 ( .A1(n5611), .A2(n5610), .A3(n5614), .ZN(n5612) );
  OAI211_X1 U6712 ( .C1(n5615), .C2(n5614), .A(n5613), .B(n5612), .ZN(n5616)
         );
  AOI21_X1 U6713 ( .B1(n6168), .B2(n5617), .A(n5616), .ZN(n5618) );
  OAI21_X1 U6714 ( .B1(n5619), .B2(n5680), .A(n5618), .ZN(U2987) );
  AOI21_X1 U6715 ( .B1(n5621), .B2(n6168), .A(n5620), .ZN(n5622) );
  OAI21_X1 U6716 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5623), .A(n5622), 
        .ZN(n5624) );
  AOI21_X1 U6717 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5625), .A(n5624), 
        .ZN(n5626) );
  OAI21_X1 U6718 ( .B1(n5627), .B2(n5680), .A(n5626), .ZN(U2989) );
  XNOR2_X1 U6719 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5633) );
  NAND3_X1 U6720 ( .A1(n5643), .A2(n5642), .A3(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5632) );
  INV_X1 U6721 ( .A(n5628), .ZN(n5630) );
  AOI21_X1 U6722 ( .B1(n5630), .B2(n6168), .A(n5629), .ZN(n5631) );
  OAI211_X1 U6723 ( .C1(n5637), .C2(n5633), .A(n5632), .B(n5631), .ZN(n5634)
         );
  AOI21_X1 U6724 ( .B1(n5635), .B2(n6171), .A(n5634), .ZN(n5636) );
  INV_X1 U6725 ( .A(n5636), .ZN(U2990) );
  INV_X1 U6726 ( .A(n5637), .ZN(n5641) );
  NOR2_X1 U6727 ( .A1(n5819), .A2(n5655), .ZN(n5639) );
  AOI211_X1 U6728 ( .C1(n5641), .C2(n5640), .A(n5639), .B(n5638), .ZN(n5645)
         );
  NAND3_X1 U6729 ( .A1(n5643), .A2(n5642), .A3(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5644) );
  OAI211_X1 U6730 ( .C1(n5646), .C2(n5680), .A(n5645), .B(n5644), .ZN(U2991)
         );
  NAND3_X1 U6731 ( .A1(n5657), .A2(n5659), .A3(n5647), .ZN(n5649) );
  OAI211_X1 U6732 ( .C1(n5655), .C2(n5838), .A(n5649), .B(n5648), .ZN(n5650)
         );
  AOI21_X1 U6733 ( .B1(n5651), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5650), 
        .ZN(n5652) );
  OAI21_X1 U6734 ( .B1(n5653), .B2(n5680), .A(n5652), .ZN(U2995) );
  OAI21_X1 U6735 ( .B1(n5656), .B2(n5655), .A(n5654), .ZN(n5661) );
  INV_X1 U6736 ( .A(n5657), .ZN(n5666) );
  NOR3_X1 U6737 ( .A1(n5666), .A2(n5659), .A3(n5658), .ZN(n5660) );
  AOI211_X1 U6738 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5668), .A(n5661), .B(n5660), .ZN(n5662) );
  OAI21_X1 U6739 ( .B1(n5663), .B2(n5680), .A(n5662), .ZN(U2996) );
  NAND2_X1 U6740 ( .A1(n5849), .A2(n6168), .ZN(n5665) );
  OAI211_X1 U6741 ( .C1(n5666), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5665), .B(n5664), .ZN(n5667) );
  AOI21_X1 U6742 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5668), .A(n5667), 
        .ZN(n5669) );
  OAI21_X1 U6743 ( .B1(n5670), .B2(n5680), .A(n5669), .ZN(U2997) );
  NAND2_X1 U6744 ( .A1(n5671), .A2(n6171), .ZN(n5677) );
  INV_X1 U6745 ( .A(n5885), .ZN(n5672) );
  NOR3_X1 U6746 ( .A1(n5672), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n5889), 
        .ZN(n5673) );
  AOI211_X1 U6747 ( .C1(n6168), .C2(n5675), .A(n5674), .B(n5673), .ZN(n5676)
         );
  OAI211_X1 U6748 ( .C1(n5679), .C2(n5678), .A(n5677), .B(n5676), .ZN(U3000)
         );
  OR2_X1 U6749 ( .A1(n5681), .A2(n5680), .ZN(n5691) );
  INV_X1 U6750 ( .A(n5682), .ZN(n5684) );
  AOI21_X1 U6751 ( .B1(n6168), .B2(n5684), .A(n5683), .ZN(n5690) );
  NAND2_X1 U6752 ( .A1(n5685), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5689)
         );
  NAND3_X1 U6753 ( .A1(n5687), .A2(n6583), .A3(n5686), .ZN(n5688) );
  NAND4_X1 U6754 ( .A1(n5691), .A2(n5690), .A3(n5689), .A4(n5688), .ZN(U3017)
         );
  OAI211_X1 U6755 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4554), .A(n6254), .B(
        n6500), .ZN(n5692) );
  OAI21_X1 U6756 ( .B1(n5694), .B2(n5693), .A(n5692), .ZN(n5695) );
  MUX2_X1 U6757 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5695), .S(n6182), 
        .Z(U3464) );
  NOR3_X1 U6758 ( .A1(n5697), .A2(n5696), .A3(n6308), .ZN(n5698) );
  AOI21_X1 U6759 ( .B1(n5699), .B2(n6222), .A(n5698), .ZN(n5700) );
  OAI21_X1 U6760 ( .B1(n6188), .B2(n5701), .A(n5700), .ZN(n5702) );
  MUX2_X1 U6761 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5702), .S(n6182), 
        .Z(U3462) );
  NOR3_X1 U6762 ( .A1(n5745), .A2(n5703), .A3(n6308), .ZN(n5705) );
  OAI21_X1 U6763 ( .B1(n5705), .B2(n6224), .A(n5704), .ZN(n5712) );
  NOR2_X1 U6764 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5706), .ZN(n5746)
         );
  INV_X1 U6765 ( .A(n5746), .ZN(n5710) );
  INV_X1 U6766 ( .A(n5755), .ZN(n5707) );
  NOR2_X1 U6767 ( .A1(n5756), .A2(n5707), .ZN(n6220) );
  OAI21_X1 U6768 ( .B1(n6220), .B2(n6405), .A(n5708), .ZN(n6225) );
  AOI211_X1 U6769 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5710), .A(n5709), .B(
        n6225), .ZN(n5711) );
  AOI22_X1 U6770 ( .A1(n5713), .A2(n6500), .B1(n6226), .B2(n6220), .ZN(n5742)
         );
  OAI22_X1 U6771 ( .A1(n5743), .A2(n6318), .B1(n5742), .B2(n5762), .ZN(n5714)
         );
  AOI21_X1 U6772 ( .B1(n5745), .B2(n6315), .A(n5714), .ZN(n5716) );
  NAND2_X1 U6773 ( .A1(n6304), .A2(n5746), .ZN(n5715) );
  OAI211_X1 U6774 ( .C1(n5750), .C2(n5717), .A(n5716), .B(n5715), .ZN(U3020)
         );
  OAI22_X1 U6775 ( .A1(n5743), .A2(n6324), .B1(n5742), .B2(n5768), .ZN(n5718)
         );
  AOI21_X1 U6776 ( .B1(n6321), .B2(n5745), .A(n5718), .ZN(n5720) );
  NAND2_X1 U6777 ( .A1(n6320), .A2(n5746), .ZN(n5719) );
  OAI211_X1 U6778 ( .C1(n5750), .C2(n5721), .A(n5720), .B(n5719), .ZN(U3021)
         );
  OAI22_X1 U6779 ( .A1(n5743), .A2(n6330), .B1(n5742), .B2(n5773), .ZN(n5722)
         );
  AOI21_X1 U6780 ( .B1(n6327), .B2(n5745), .A(n5722), .ZN(n5724) );
  NAND2_X1 U6781 ( .A1(n6326), .A2(n5746), .ZN(n5723) );
  OAI211_X1 U6782 ( .C1(n5750), .C2(n5725), .A(n5724), .B(n5723), .ZN(U3022)
         );
  INV_X1 U6783 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5729) );
  OAI22_X1 U6784 ( .A1(n5743), .A2(n6336), .B1(n5742), .B2(n5778), .ZN(n5726)
         );
  AOI21_X1 U6785 ( .B1(n6333), .B2(n5745), .A(n5726), .ZN(n5728) );
  NAND2_X1 U6786 ( .A1(n6332), .A2(n5746), .ZN(n5727) );
  OAI211_X1 U6787 ( .C1(n5750), .C2(n5729), .A(n5728), .B(n5727), .ZN(U3023)
         );
  OAI22_X1 U6788 ( .A1(n5743), .A2(n6342), .B1(n5742), .B2(n5783), .ZN(n5730)
         );
  AOI21_X1 U6789 ( .B1(n6339), .B2(n5745), .A(n5730), .ZN(n5732) );
  NAND2_X1 U6790 ( .A1(n6338), .A2(n5746), .ZN(n5731) );
  OAI211_X1 U6791 ( .C1(n5750), .C2(n5733), .A(n5732), .B(n5731), .ZN(U3024)
         );
  OAI22_X1 U6792 ( .A1(n5743), .A2(n6348), .B1(n5742), .B2(n5788), .ZN(n5734)
         );
  AOI21_X1 U6793 ( .B1(n6345), .B2(n5745), .A(n5734), .ZN(n5736) );
  NAND2_X1 U6794 ( .A1(n6344), .A2(n5746), .ZN(n5735) );
  OAI211_X1 U6795 ( .C1(n5750), .C2(n5737), .A(n5736), .B(n5735), .ZN(U3025)
         );
  OAI22_X1 U6796 ( .A1(n5743), .A2(n6354), .B1(n5742), .B2(n5793), .ZN(n5738)
         );
  AOI21_X1 U6797 ( .B1(n6351), .B2(n5745), .A(n5738), .ZN(n5740) );
  NAND2_X1 U6798 ( .A1(n6350), .A2(n5746), .ZN(n5739) );
  OAI211_X1 U6799 ( .C1(n5750), .C2(n5741), .A(n5740), .B(n5739), .ZN(U3026)
         );
  OAI22_X1 U6800 ( .A1(n5743), .A2(n6365), .B1(n5742), .B2(n5798), .ZN(n5744)
         );
  AOI21_X1 U6801 ( .B1(n6360), .B2(n5745), .A(n5744), .ZN(n5748) );
  NAND2_X1 U6802 ( .A1(n6358), .A2(n5746), .ZN(n5747) );
  OAI211_X1 U6803 ( .C1(n5750), .C2(n5749), .A(n5748), .B(n5747), .ZN(U3027)
         );
  NAND3_X1 U6804 ( .A1(n5801), .A2(n6500), .A3(n5800), .ZN(n5753) );
  NOR2_X1 U6805 ( .A1(n6301), .A2(n5751), .ZN(n5761) );
  AOI21_X1 U6806 ( .B1(n5753), .B2(n5752), .A(n5761), .ZN(n5759) );
  NOR2_X1 U6807 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5754), .ZN(n5804)
         );
  OR2_X1 U6808 ( .A1(n5756), .A2(n5755), .ZN(n6299) );
  AOI21_X1 U6809 ( .B1(n6299), .B2(STATE2_REG_2__SCAN_IN), .A(n5757), .ZN(
        n6311) );
  OAI211_X1 U6810 ( .C1(n6483), .C2(n5804), .A(n6300), .B(n6311), .ZN(n5758)
         );
  INV_X1 U6811 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5767) );
  INV_X1 U6812 ( .A(n6299), .ZN(n5760) );
  AOI22_X1 U6813 ( .A1(n5761), .A2(n6500), .B1(n6226), .B2(n5760), .ZN(n5799)
         );
  OAI22_X1 U6814 ( .A1(n5800), .A2(n6318), .B1(n5799), .B2(n5762), .ZN(n5763)
         );
  AOI21_X1 U6815 ( .B1(n5764), .B2(n6315), .A(n5763), .ZN(n5766) );
  NAND2_X1 U6816 ( .A1(n6304), .A2(n5804), .ZN(n5765) );
  OAI211_X1 U6817 ( .C1(n5807), .C2(n5767), .A(n5766), .B(n5765), .ZN(U3084)
         );
  INV_X1 U6818 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5772) );
  OAI22_X1 U6819 ( .A1(n5800), .A2(n6324), .B1(n5799), .B2(n5768), .ZN(n5770)
         );
  NOR2_X1 U6820 ( .A1(n5801), .A2(n6269), .ZN(n5769) );
  AOI211_X1 U6821 ( .C1(n5804), .C2(n6320), .A(n5770), .B(n5769), .ZN(n5771)
         );
  OAI21_X1 U6822 ( .B1(n5807), .B2(n5772), .A(n5771), .ZN(U3085) );
  INV_X1 U6823 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5777) );
  OAI22_X1 U6824 ( .A1(n5800), .A2(n6330), .B1(n5799), .B2(n5773), .ZN(n5775)
         );
  NOR2_X1 U6825 ( .A1(n5801), .A2(n6273), .ZN(n5774) );
  AOI211_X1 U6826 ( .C1(n5804), .C2(n6326), .A(n5775), .B(n5774), .ZN(n5776)
         );
  OAI21_X1 U6827 ( .B1(n5807), .B2(n5777), .A(n5776), .ZN(U3086) );
  INV_X1 U6828 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5782) );
  OAI22_X1 U6829 ( .A1(n5800), .A2(n6336), .B1(n5799), .B2(n5778), .ZN(n5780)
         );
  NOR2_X1 U6830 ( .A1(n5801), .A2(n6277), .ZN(n5779) );
  AOI211_X1 U6831 ( .C1(n5804), .C2(n6332), .A(n5780), .B(n5779), .ZN(n5781)
         );
  OAI21_X1 U6832 ( .B1(n5807), .B2(n5782), .A(n5781), .ZN(U3087) );
  INV_X1 U6833 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5787) );
  OAI22_X1 U6834 ( .A1(n5800), .A2(n6342), .B1(n5799), .B2(n5783), .ZN(n5785)
         );
  NOR2_X1 U6835 ( .A1(n5801), .A2(n6281), .ZN(n5784) );
  AOI211_X1 U6836 ( .C1(n5804), .C2(n6338), .A(n5785), .B(n5784), .ZN(n5786)
         );
  OAI21_X1 U6837 ( .B1(n5807), .B2(n5787), .A(n5786), .ZN(U3088) );
  INV_X1 U6838 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5792) );
  OAI22_X1 U6839 ( .A1(n5800), .A2(n6348), .B1(n5799), .B2(n5788), .ZN(n5790)
         );
  NOR2_X1 U6840 ( .A1(n5801), .A2(n6285), .ZN(n5789) );
  AOI211_X1 U6841 ( .C1(n5804), .C2(n6344), .A(n5790), .B(n5789), .ZN(n5791)
         );
  OAI21_X1 U6842 ( .B1(n5807), .B2(n5792), .A(n5791), .ZN(U3089) );
  INV_X1 U6843 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5797) );
  OAI22_X1 U6844 ( .A1(n5800), .A2(n6354), .B1(n5799), .B2(n5793), .ZN(n5795)
         );
  NOR2_X1 U6845 ( .A1(n5801), .A2(n6290), .ZN(n5794) );
  AOI211_X1 U6846 ( .C1(n5804), .C2(n6350), .A(n5795), .B(n5794), .ZN(n5796)
         );
  OAI21_X1 U6847 ( .B1(n5807), .B2(n5797), .A(n5796), .ZN(U3090) );
  INV_X1 U6848 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5806) );
  OAI22_X1 U6849 ( .A1(n5800), .A2(n6365), .B1(n5799), .B2(n5798), .ZN(n5803)
         );
  NOR2_X1 U6850 ( .A1(n5801), .A2(n6218), .ZN(n5802) );
  AOI211_X1 U6851 ( .C1(n5804), .C2(n6358), .A(n5803), .B(n5802), .ZN(n5805)
         );
  OAI21_X1 U6852 ( .B1(n5807), .B2(n5806), .A(n5805), .ZN(U3091) );
  AND2_X1 U6853 ( .A1(n6032), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U6854 ( .A(n5808), .ZN(n5809) );
  AOI21_X1 U6855 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n5810), .A(n5809), .ZN(
        n5811) );
  NAND2_X1 U6856 ( .A1(n5812), .A2(n5811), .ZN(U2788) );
  OAI22_X1 U6857 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5814), .B1(n5813), .B2(
        n5997), .ZN(n5818) );
  OAI22_X1 U6858 ( .A1(n5816), .A2(n6464), .B1(n3852), .B2(n5815), .ZN(n5817)
         );
  AOI211_X1 U6859 ( .C1(EBX_REG_27__SCAN_IN), .C2(n5993), .A(n5818), .B(n5817), 
        .ZN(n5824) );
  OAI22_X1 U6860 ( .A1(n5821), .A2(n5820), .B1(n5819), .B2(n5983), .ZN(n5822)
         );
  INV_X1 U6861 ( .A(n5822), .ZN(n5823) );
  NAND2_X1 U6862 ( .A1(n5824), .A2(n5823), .ZN(U2800) );
  INV_X1 U6863 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6462) );
  AOI22_X1 U6864 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n5991), .B1(n5825), 
        .B2(n6462), .ZN(n5835) );
  AOI22_X1 U6865 ( .A1(EBX_REG_25__SCAN_IN), .A2(n5993), .B1(n5826), .B2(n5958), .ZN(n5834) );
  NOR2_X1 U6866 ( .A1(n5827), .A2(n5983), .ZN(n5828) );
  AOI21_X1 U6867 ( .B1(n5829), .B2(n5976), .A(n5828), .ZN(n5833) );
  INV_X1 U6868 ( .A(n5839), .ZN(n5830) );
  OAI21_X1 U6869 ( .B1(n5831), .B2(n5830), .A(REIP_REG_25__SCAN_IN), .ZN(n5832) );
  NAND4_X1 U6870 ( .A1(n5835), .A2(n5834), .A3(n5833), .A4(n5832), .ZN(U2802)
         );
  AOI22_X1 U6871 ( .A1(EBX_REG_23__SCAN_IN), .A2(n5993), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n5991), .ZN(n5843) );
  AOI21_X1 U6872 ( .B1(n5837), .B2(n5836), .A(REIP_REG_23__SCAN_IN), .ZN(n5840) );
  OAI22_X1 U6873 ( .A1(n5840), .A2(n5839), .B1(n5838), .B2(n5983), .ZN(n5841)
         );
  AOI21_X1 U6874 ( .B1(n5863), .B2(n5976), .A(n5841), .ZN(n5842) );
  OAI211_X1 U6875 ( .C1(n5844), .C2(n5997), .A(n5843), .B(n5842), .ZN(U2804)
         );
  AOI22_X1 U6876 ( .A1(EBX_REG_21__SCAN_IN), .A2(n5993), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n5991), .ZN(n5845) );
  OAI221_X1 U6877 ( .B1(n5847), .B2(n6457), .C1(n5846), .C2(
        REIP_REG_21__SCAN_IN), .A(n5845), .ZN(n5848) );
  INV_X1 U6878 ( .A(n5848), .ZN(n5851) );
  AOI22_X1 U6879 ( .A1(n5866), .A2(n5976), .B1(n5992), .B2(n5849), .ZN(n5850)
         );
  OAI211_X1 U6880 ( .C1(n5852), .C2(n5997), .A(n5851), .B(n5850), .ZN(U2806)
         );
  AOI211_X1 U6881 ( .C1(n5084), .C2(n6453), .A(n5854), .B(n5853), .ZN(n5855)
         );
  AOI211_X1 U6882 ( .C1(n5991), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5855), 
        .B(n5956), .ZN(n5856) );
  OAI21_X1 U6883 ( .B1(n5084), .B2(n5931), .A(n5856), .ZN(n5857) );
  AOI21_X1 U6884 ( .B1(EBX_REG_19__SCAN_IN), .B2(n5993), .A(n5857), .ZN(n5860)
         );
  AOI22_X1 U6885 ( .A1(n5872), .A2(n5976), .B1(n5992), .B2(n5858), .ZN(n5859)
         );
  OAI211_X1 U6886 ( .C1(n5861), .C2(n5997), .A(n5860), .B(n5859), .ZN(U2808)
         );
  INV_X1 U6887 ( .A(n5862), .ZN(n6012) );
  AOI22_X1 U6888 ( .A1(n5863), .A2(n6012), .B1(n6011), .B2(DATAI_7_), .ZN(
        n5865) );
  AOI22_X1 U6889 ( .A1(n6015), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6014), .ZN(n5864) );
  NAND2_X1 U6890 ( .A1(n5865), .A2(n5864), .ZN(U2868) );
  AOI22_X1 U6891 ( .A1(n5866), .A2(n6012), .B1(n6011), .B2(DATAI_5_), .ZN(
        n5868) );
  AOI22_X1 U6892 ( .A1(n6015), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n6014), .ZN(n5867) );
  NAND2_X1 U6893 ( .A1(n5868), .A2(n5867), .ZN(U2870) );
  AOI22_X1 U6894 ( .A1(n5869), .A2(n6012), .B1(n6011), .B2(DATAI_4_), .ZN(
        n5871) );
  AOI22_X1 U6895 ( .A1(n6015), .A2(DATAI_20_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n6014), .ZN(n5870) );
  NAND2_X1 U6896 ( .A1(n5871), .A2(n5870), .ZN(U2871) );
  AOI22_X1 U6897 ( .A1(n5872), .A2(n6012), .B1(n6011), .B2(DATAI_3_), .ZN(
        n5874) );
  AOI22_X1 U6898 ( .A1(n6015), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6014), .ZN(n5873) );
  NAND2_X1 U6899 ( .A1(n5874), .A2(n5873), .ZN(U2872) );
  AOI22_X1 U6900 ( .A1(n6167), .A2(REIP_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6109), .ZN(n5884) );
  INV_X1 U6901 ( .A(n5876), .ZN(n5878) );
  NAND3_X1 U6902 ( .A1(n5876), .A2(n5875), .A3(n5579), .ZN(n5877) );
  AOI22_X1 U6903 ( .A1(n5878), .A2(n5581), .B1(n5877), .B2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5882) );
  INV_X1 U6904 ( .A(n5879), .ZN(n5880) );
  OAI21_X1 U6905 ( .B1(n5882), .B2(n5881), .A(n5880), .ZN(n5886) );
  AOI22_X1 U6906 ( .A1(n5886), .A2(n6114), .B1(n2946), .B2(n6008), .ZN(n5883)
         );
  OAI211_X1 U6907 ( .C1(n5937), .C2(n6118), .A(n5884), .B(n5883), .ZN(U2969)
         );
  AOI22_X1 U6908 ( .A1(n6167), .A2(REIP_REG_17__SCAN_IN), .B1(n5889), .B2(
        n5885), .ZN(n5888) );
  AOI22_X1 U6909 ( .A1(n5886), .A2(n6171), .B1(n6168), .B2(n5934), .ZN(n5887)
         );
  OAI211_X1 U6910 ( .C1(n5890), .C2(n5889), .A(n5888), .B(n5887), .ZN(U3001)
         );
  INV_X1 U6911 ( .A(n5945), .ZN(n5892) );
  AOI21_X1 U6912 ( .B1(n6168), .B2(n5892), .A(n5891), .ZN(n5896) );
  AOI22_X1 U6913 ( .A1(n5894), .A2(n6171), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5893), .ZN(n5895) );
  OAI211_X1 U6914 ( .C1(n5898), .C2(n5897), .A(n5896), .B(n5895), .ZN(U3005)
         );
  NAND4_X1 U6915 ( .A1(n5902), .A2(n5901), .A3(n5900), .A4(n5899), .ZN(n5903)
         );
  OAI21_X1 U6916 ( .B1(n5904), .B2(n6607), .A(n5903), .ZN(U3455) );
  AOI21_X1 U6917 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6548), .A(n6424), .ZN(n5910) );
  INV_X1 U6918 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5905) );
  AND2_X1 U6919 ( .A1(STATE_REG_1__SCAN_IN), .A2(n6424), .ZN(n6512) );
  AOI21_X1 U6920 ( .B1(n5910), .B2(n5905), .A(n6512), .ZN(U2789) );
  INV_X1 U6921 ( .A(n5906), .ZN(n5907) );
  OAI21_X1 U6922 ( .B1(n5907), .B2(n6407), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5908) );
  OAI21_X1 U6923 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6408), .A(n5908), .ZN(
        U2790) );
  INV_X1 U6924 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6532) );
  NOR2_X1 U6925 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5911) );
  NOR2_X1 U6926 ( .A1(n6512), .A2(n5911), .ZN(n5909) );
  AOI22_X1 U6927 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n6512), .B1(n6532), .B2(
        n5909), .ZN(U2791) );
  NOR2_X1 U6928 ( .A1(n6512), .A2(n5910), .ZN(n6479) );
  OAI21_X1 U6929 ( .B1(BS16_N), .B2(n5911), .A(n6479), .ZN(n6477) );
  OAI21_X1 U6930 ( .B1(n6479), .B2(n6305), .A(n6477), .ZN(U2792) );
  OAI21_X1 U6931 ( .B1(n5914), .B2(n5913), .A(n5912), .ZN(U2793) );
  NOR4_X1 U6932 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n5918) );
  NOR4_X1 U6933 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n5917) );
  NOR4_X1 U6934 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5916) );
  NOR4_X1 U6935 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n5915) );
  NAND4_X1 U6936 ( .A1(n5918), .A2(n5917), .A3(n5916), .A4(n5915), .ZN(n5924)
         );
  NOR4_X1 U6937 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_26__SCAN_IN), .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n5922) );
  AOI211_X1 U6938 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_16__SCAN_IN), .B(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n5921) );
  NOR4_X1 U6939 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n5920) );
  NOR4_X1 U6940 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n5919) );
  NAND4_X1 U6941 ( .A1(n5922), .A2(n5921), .A3(n5920), .A4(n5919), .ZN(n5923)
         );
  NOR2_X1 U6942 ( .A1(n5924), .A2(n5923), .ZN(n6497) );
  INV_X1 U6943 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5926) );
  NOR3_X1 U6944 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5927) );
  OAI21_X1 U6945 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5927), .A(n6497), .ZN(n5925)
         );
  OAI21_X1 U6946 ( .B1(n6497), .B2(n5926), .A(n5925), .ZN(U2794) );
  INV_X1 U6947 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6478) );
  AOI21_X1 U6948 ( .B1(n6490), .B2(n6478), .A(n5927), .ZN(n5929) );
  INV_X1 U6949 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5928) );
  INV_X1 U6950 ( .A(n6497), .ZN(n6492) );
  AOI22_X1 U6951 ( .A1(n6497), .A2(n5929), .B1(n5928), .B2(n6492), .ZN(U2795)
         );
  AOI21_X1 U6952 ( .B1(REIP_REG_16__SCAN_IN), .B2(n5930), .A(
        REIP_REG_17__SCAN_IN), .ZN(n5932) );
  OAI22_X1 U6953 ( .A1(n5932), .A2(n5931), .B1(n6623), .B2(n5954), .ZN(n5933)
         );
  AOI211_X1 U6954 ( .C1(n5991), .C2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n5956), 
        .B(n5933), .ZN(n5936) );
  AOI22_X1 U6955 ( .A1(n6008), .A2(n5976), .B1(n5992), .B2(n5934), .ZN(n5935)
         );
  OAI211_X1 U6956 ( .C1(n5937), .C2(n5997), .A(n5936), .B(n5935), .ZN(U2810)
         );
  INV_X1 U6957 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6445) );
  AOI21_X1 U6958 ( .B1(n5939), .B2(n6445), .A(n5938), .ZN(n5952) );
  NAND2_X1 U6959 ( .A1(n5991), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5940)
         );
  OAI211_X1 U6960 ( .C1(REIP_REG_13__SCAN_IN), .C2(n5941), .A(n5940), .B(n5982), .ZN(n5942) );
  INV_X1 U6961 ( .A(n5942), .ZN(n5944) );
  NAND2_X1 U6962 ( .A1(n5993), .A2(EBX_REG_13__SCAN_IN), .ZN(n5943) );
  OAI211_X1 U6963 ( .C1(n5945), .C2(n5983), .A(n5944), .B(n5943), .ZN(n5946)
         );
  INV_X1 U6964 ( .A(n5946), .ZN(n5951) );
  INV_X1 U6965 ( .A(n5947), .ZN(n5948) );
  AOI22_X1 U6966 ( .A1(n5949), .A2(n5976), .B1(n5948), .B2(n5958), .ZN(n5950)
         );
  OAI211_X1 U6967 ( .C1(n5952), .C2(n5122), .A(n5951), .B(n5950), .ZN(U2814)
         );
  OAI22_X1 U6968 ( .A1(n5954), .A2(n3036), .B1(n5983), .B2(n5953), .ZN(n5955)
         );
  AOI211_X1 U6969 ( .C1(n5991), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5956), 
        .B(n5955), .ZN(n5966) );
  AOI22_X1 U6970 ( .A1(n5959), .A2(n5976), .B1(n5958), .B2(n5957), .ZN(n5965)
         );
  OAI21_X1 U6971 ( .B1(n5961), .B2(n5960), .A(REIP_REG_10__SCAN_IN), .ZN(n5964) );
  NAND3_X1 U6972 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5962), .A3(n6442), .ZN(n5963) );
  NAND4_X1 U6973 ( .A1(n5966), .A2(n5965), .A3(n5964), .A4(n5963), .ZN(U2817)
         );
  OAI21_X1 U6974 ( .B1(REIP_REG_7__SCAN_IN), .B2(REIP_REG_6__SCAN_IN), .A(
        n5967), .ZN(n5974) );
  INV_X1 U6975 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6554) );
  OR2_X1 U6976 ( .A1(n5986), .A2(n6554), .ZN(n5972) );
  NAND2_X1 U6977 ( .A1(n5993), .A2(EBX_REG_7__SCAN_IN), .ZN(n5970) );
  OR2_X1 U6978 ( .A1(n5983), .A2(n6135), .ZN(n5969) );
  NAND2_X1 U6979 ( .A1(n5991), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5968)
         );
  AND4_X1 U6980 ( .A1(n5970), .A2(n5982), .A3(n5969), .A4(n5968), .ZN(n5971)
         );
  OAI211_X1 U6981 ( .C1(n5974), .C2(n5973), .A(n5972), .B(n5971), .ZN(n5975)
         );
  AOI21_X1 U6982 ( .B1(n5976), .B2(n6089), .A(n5975), .ZN(n5977) );
  OAI21_X1 U6983 ( .B1(n6092), .B2(n5997), .A(n5977), .ZN(U2820) );
  INV_X1 U6984 ( .A(n5978), .ZN(n5980) );
  AOI21_X1 U6985 ( .B1(n5980), .B2(n5979), .A(REIP_REG_5__SCAN_IN), .ZN(n5987)
         );
  NAND2_X1 U6986 ( .A1(n5991), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5981)
         );
  OAI211_X1 U6987 ( .C1(n5983), .C2(n6145), .A(n5982), .B(n5981), .ZN(n5984)
         );
  AOI21_X1 U6988 ( .B1(n5993), .B2(EBX_REG_5__SCAN_IN), .A(n5984), .ZN(n5985)
         );
  OAI21_X1 U6989 ( .B1(n5987), .B2(n5986), .A(n5985), .ZN(n5988) );
  AOI21_X1 U6990 ( .B1(n6000), .B2(n6097), .A(n5988), .ZN(n5989) );
  OAI21_X1 U6991 ( .B1(n6100), .B2(n5997), .A(n5989), .ZN(U2822) );
  INV_X1 U6992 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U6993 ( .A1(n5990), .A2(REIP_REG_2__SCAN_IN), .ZN(n6002) );
  AOI22_X1 U6994 ( .A1(n5992), .A2(n6160), .B1(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .B2(n5991), .ZN(n5995) );
  NAND2_X1 U6995 ( .A1(n5993), .A2(EBX_REG_3__SCAN_IN), .ZN(n5994) );
  OAI211_X1 U6996 ( .C1(n6301), .C2(n5996), .A(n5995), .B(n5994), .ZN(n5999)
         );
  NOR2_X1 U6997 ( .A1(n5997), .A2(n6108), .ZN(n5998) );
  AOI211_X1 U6998 ( .C1(n6105), .C2(n6000), .A(n5999), .B(n5998), .ZN(n6001)
         );
  OAI221_X1 U6999 ( .B1(n6003), .B2(n6529), .C1(n6003), .C2(n6002), .A(n6001), 
        .ZN(U2824) );
  INV_X1 U7000 ( .A(n6004), .ZN(n6005) );
  AOI22_X1 U7001 ( .A1(n6005), .A2(n6012), .B1(n6011), .B2(DATAI_2_), .ZN(
        n6007) );
  AOI22_X1 U7002 ( .A1(n6015), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n6014), .ZN(n6006) );
  NAND2_X1 U7003 ( .A1(n6007), .A2(n6006), .ZN(U2873) );
  AOI22_X1 U7004 ( .A1(n6008), .A2(n6012), .B1(n6011), .B2(DATAI_1_), .ZN(
        n6010) );
  AOI22_X1 U7005 ( .A1(n6015), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n6014), .ZN(n6009) );
  NAND2_X1 U7006 ( .A1(n6010), .A2(n6009), .ZN(U2874) );
  AOI22_X1 U7007 ( .A1(n6013), .A2(n6012), .B1(n6011), .B2(DATAI_0_), .ZN(
        n6017) );
  AOI22_X1 U7008 ( .A1(n6015), .A2(DATAI_16_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n6014), .ZN(n6016) );
  NAND2_X1 U7009 ( .A1(n6017), .A2(n6016), .ZN(U2875) );
  INV_X1 U7010 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n6614) );
  AOI22_X1 U7011 ( .A1(EAX_REG_15__SCAN_IN), .A2(n6020), .B1(n6032), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6018) );
  OAI21_X1 U7012 ( .B1(n6395), .B2(n6614), .A(n6018), .ZN(U2908) );
  INV_X1 U7013 ( .A(LWORD_REG_14__SCAN_IN), .ZN(n6561) );
  AOI22_X1 U7014 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6020), .B1(n6032), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6019) );
  OAI21_X1 U7015 ( .B1(n6395), .B2(n6561), .A(n6019), .ZN(U2909) );
  AOI22_X1 U7016 ( .A1(n6041), .A2(LWORD_REG_13__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6021) );
  OAI21_X1 U7017 ( .B1(n6022), .B2(n6043), .A(n6021), .ZN(U2910) );
  INV_X1 U7018 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6076) );
  AOI22_X1 U7019 ( .A1(n6041), .A2(LWORD_REG_12__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6023) );
  OAI21_X1 U7020 ( .B1(n6076), .B2(n6043), .A(n6023), .ZN(U2911) );
  INV_X1 U7021 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6071) );
  AOI22_X1 U7022 ( .A1(n6041), .A2(LWORD_REG_11__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6024) );
  OAI21_X1 U7023 ( .B1(n6071), .B2(n6043), .A(n6024), .ZN(U2912) );
  INV_X1 U7024 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6068) );
  AOI22_X1 U7025 ( .A1(n6041), .A2(LWORD_REG_10__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6025) );
  OAI21_X1 U7026 ( .B1(n6068), .B2(n6043), .A(n6025), .ZN(U2913) );
  INV_X1 U7027 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6065) );
  AOI22_X1 U7028 ( .A1(n6041), .A2(LWORD_REG_9__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6026) );
  OAI21_X1 U7029 ( .B1(n6065), .B2(n6043), .A(n6026), .ZN(U2914) );
  INV_X1 U7030 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6062) );
  AOI22_X1 U7031 ( .A1(n6041), .A2(LWORD_REG_8__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6027) );
  OAI21_X1 U7032 ( .B1(n6062), .B2(n6043), .A(n6027), .ZN(U2915) );
  AOI22_X1 U7033 ( .A1(n6041), .A2(LWORD_REG_7__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6028) );
  OAI21_X1 U7034 ( .B1(n6029), .B2(n6043), .A(n6028), .ZN(U2916) );
  AOI22_X1 U7035 ( .A1(n6501), .A2(LWORD_REG_6__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6030) );
  OAI21_X1 U7036 ( .B1(n6537), .B2(n6043), .A(n6030), .ZN(U2917) );
  AOI22_X1 U7037 ( .A1(n6501), .A2(LWORD_REG_5__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6031) );
  OAI21_X1 U7038 ( .B1(n4309), .B2(n6043), .A(n6031), .ZN(U2918) );
  AOI22_X1 U7039 ( .A1(n6501), .A2(LWORD_REG_4__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6033) );
  OAI21_X1 U7040 ( .B1(n6034), .B2(n6043), .A(n6033), .ZN(U2919) );
  INV_X1 U7041 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6586) );
  AOI22_X1 U7042 ( .A1(n6501), .A2(LWORD_REG_3__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6035) );
  OAI21_X1 U7043 ( .B1(n6586), .B2(n6043), .A(n6035), .ZN(U2920) );
  AOI22_X1 U7044 ( .A1(n6501), .A2(LWORD_REG_2__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6036) );
  OAI21_X1 U7045 ( .B1(n6037), .B2(n6043), .A(n6036), .ZN(U2921) );
  AOI22_X1 U7046 ( .A1(n6501), .A2(LWORD_REG_1__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6038) );
  OAI21_X1 U7047 ( .B1(n6039), .B2(n6043), .A(n6038), .ZN(U2922) );
  AOI22_X1 U7048 ( .A1(n6041), .A2(LWORD_REG_0__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6042) );
  OAI21_X1 U7049 ( .B1(n6044), .B2(n6043), .A(n6042), .ZN(U2923) );
  INV_X1 U7050 ( .A(DATAI_8_), .ZN(n6045) );
  NOR2_X1 U7051 ( .A1(n6058), .A2(n6045), .ZN(n6060) );
  AOI21_X1 U7052 ( .B1(n6073), .B2(UWORD_REG_8__SCAN_IN), .A(n6060), .ZN(n6046) );
  OAI21_X1 U7053 ( .B1(n6047), .B2(n6075), .A(n6046), .ZN(U2932) );
  INV_X1 U7054 ( .A(DATAI_9_), .ZN(n6048) );
  NOR2_X1 U7055 ( .A1(n6058), .A2(n6048), .ZN(n6063) );
  AOI21_X1 U7056 ( .B1(n6073), .B2(UWORD_REG_9__SCAN_IN), .A(n6063), .ZN(n6049) );
  OAI21_X1 U7057 ( .B1(n6050), .B2(n6075), .A(n6049), .ZN(U2933) );
  INV_X1 U7058 ( .A(DATAI_10_), .ZN(n6051) );
  NOR2_X1 U7059 ( .A1(n6058), .A2(n6051), .ZN(n6066) );
  AOI21_X1 U7060 ( .B1(n6073), .B2(UWORD_REG_10__SCAN_IN), .A(n6066), .ZN(
        n6052) );
  OAI21_X1 U7061 ( .B1(n3866), .B2(n6075), .A(n6052), .ZN(U2934) );
  INV_X1 U7062 ( .A(DATAI_11_), .ZN(n6053) );
  NOR2_X1 U7063 ( .A1(n6058), .A2(n6053), .ZN(n6069) );
  AOI21_X1 U7064 ( .B1(n6073), .B2(UWORD_REG_11__SCAN_IN), .A(n6069), .ZN(
        n6054) );
  OAI21_X1 U7065 ( .B1(n3859), .B2(n6075), .A(n6054), .ZN(U2935) );
  INV_X1 U7066 ( .A(DATAI_12_), .ZN(n6055) );
  NOR2_X1 U7067 ( .A1(n6058), .A2(n6055), .ZN(n6072) );
  AOI21_X1 U7068 ( .B1(n6073), .B2(UWORD_REG_12__SCAN_IN), .A(n6072), .ZN(
        n6056) );
  OAI21_X1 U7069 ( .B1(n6609), .B2(n6075), .A(n6056), .ZN(U2936) );
  INV_X1 U7070 ( .A(DATAI_14_), .ZN(n6057) );
  NOR2_X1 U7071 ( .A1(n6058), .A2(n6057), .ZN(n6077) );
  AOI21_X1 U7072 ( .B1(n6073), .B2(UWORD_REG_14__SCAN_IN), .A(n6077), .ZN(
        n6059) );
  OAI21_X1 U7073 ( .B1(n3955), .B2(n6075), .A(n6059), .ZN(U2938) );
  AOI21_X1 U7074 ( .B1(n6073), .B2(LWORD_REG_8__SCAN_IN), .A(n6060), .ZN(n6061) );
  OAI21_X1 U7075 ( .B1(n6062), .B2(n6075), .A(n6061), .ZN(U2947) );
  AOI21_X1 U7076 ( .B1(n6073), .B2(LWORD_REG_9__SCAN_IN), .A(n6063), .ZN(n6064) );
  OAI21_X1 U7077 ( .B1(n6065), .B2(n6075), .A(n6064), .ZN(U2948) );
  AOI21_X1 U7078 ( .B1(n6073), .B2(LWORD_REG_10__SCAN_IN), .A(n6066), .ZN(
        n6067) );
  OAI21_X1 U7079 ( .B1(n6068), .B2(n6075), .A(n6067), .ZN(U2949) );
  AOI21_X1 U7080 ( .B1(n6073), .B2(LWORD_REG_11__SCAN_IN), .A(n6069), .ZN(
        n6070) );
  OAI21_X1 U7081 ( .B1(n6071), .B2(n6075), .A(n6070), .ZN(U2950) );
  AOI21_X1 U7082 ( .B1(n6073), .B2(LWORD_REG_12__SCAN_IN), .A(n6072), .ZN(
        n6074) );
  OAI21_X1 U7083 ( .B1(n6076), .B2(n6075), .A(n6074), .ZN(U2951) );
  AOI21_X1 U7084 ( .B1(n6079), .B2(EAX_REG_14__SCAN_IN), .A(n6077), .ZN(n6078)
         );
  OAI21_X1 U7085 ( .B1(n6561), .B2(n6082), .A(n6078), .ZN(U2953) );
  AOI22_X1 U7086 ( .A1(n6080), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6079), .ZN(n6081) );
  OAI21_X1 U7087 ( .B1(n6614), .B2(n6082), .A(n6081), .ZN(U2954) );
  AOI22_X1 U7088 ( .A1(n6167), .A2(REIP_REG_7__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n6109), .ZN(n6091) );
  NAND2_X1 U7089 ( .A1(n6084), .A2(n6083), .ZN(n6087) );
  OAI21_X1 U7090 ( .B1(n6087), .B2(n6086), .A(n6085), .ZN(n6088) );
  INV_X1 U7091 ( .A(n6088), .ZN(n6138) );
  AOI22_X1 U7092 ( .A1(n6138), .A2(n6114), .B1(n2946), .B2(n6089), .ZN(n6090)
         );
  OAI211_X1 U7093 ( .C1(n6092), .C2(n6118), .A(n6091), .B(n6090), .ZN(U2979)
         );
  AOI22_X1 U7094 ( .A1(n6167), .A2(REIP_REG_5__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n6109), .ZN(n6099) );
  OAI21_X1 U7095 ( .B1(n6095), .B2(n6094), .A(n6093), .ZN(n6096) );
  INV_X1 U7096 ( .A(n6096), .ZN(n6147) );
  AOI22_X1 U7097 ( .A1(n6147), .A2(n6114), .B1(n2946), .B2(n6097), .ZN(n6098)
         );
  OAI211_X1 U7098 ( .C1(n6100), .C2(n6118), .A(n6099), .B(n6098), .ZN(U2981)
         );
  AOI22_X1 U7099 ( .A1(n6167), .A2(REIP_REG_3__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n6109), .ZN(n6107) );
  OR2_X1 U7100 ( .A1(n6102), .A2(n6101), .ZN(n6104) );
  AND2_X1 U7101 ( .A1(n6104), .A2(n6103), .ZN(n6161) );
  AOI22_X1 U7102 ( .A1(n6114), .A2(n6161), .B1(n6105), .B2(n2946), .ZN(n6106)
         );
  OAI211_X1 U7103 ( .C1(n6108), .C2(n6118), .A(n6107), .B(n6106), .ZN(U2983)
         );
  AOI22_X1 U7104 ( .A1(n6167), .A2(REIP_REG_2__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6109), .ZN(n6117) );
  INV_X1 U7105 ( .A(n6110), .ZN(n6115) );
  XOR2_X1 U7106 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .B(n6111), .Z(n6113) );
  XNOR2_X1 U7107 ( .A(n6113), .B(n6112), .ZN(n6170) );
  AOI22_X1 U7108 ( .A1(n6115), .A2(n2946), .B1(n6114), .B2(n6170), .ZN(n6116)
         );
  OAI211_X1 U7109 ( .C1(n6119), .C2(n6118), .A(n6117), .B(n6116), .ZN(U2984)
         );
  AOI21_X1 U7110 ( .B1(n6168), .B2(n6121), .A(n6120), .ZN(n6125) );
  AOI22_X1 U7111 ( .A1(n6171), .A2(n6123), .B1(n6126), .B2(n6122), .ZN(n6124)
         );
  OAI211_X1 U7112 ( .C1(n6127), .C2(n6126), .A(n6125), .B(n6124), .ZN(U3007)
         );
  AOI21_X1 U7113 ( .B1(n6168), .B2(n6129), .A(n6128), .ZN(n6133) );
  AOI22_X1 U7114 ( .A1(n6131), .A2(n6171), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6130), .ZN(n6132) );
  OAI211_X1 U7115 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6134), .A(n6133), 
        .B(n6132), .ZN(U3009) );
  INV_X1 U7116 ( .A(n6135), .ZN(n6136) );
  AOI22_X1 U7117 ( .A1(n6168), .A2(n6136), .B1(n6167), .B2(REIP_REG_7__SCAN_IN), .ZN(n6140) );
  AOI22_X1 U7118 ( .A1(n6138), .A2(n6171), .B1(n6137), .B2(n6141), .ZN(n6139)
         );
  OAI211_X1 U7119 ( .C1(n6142), .C2(n6141), .A(n6140), .B(n6139), .ZN(U3011)
         );
  INV_X1 U7120 ( .A(n6155), .ZN(n6143) );
  AOI21_X1 U7121 ( .B1(n6144), .B2(n6143), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6150) );
  INV_X1 U7122 ( .A(n6145), .ZN(n6146) );
  AOI22_X1 U7123 ( .A1(n6147), .A2(n6171), .B1(n6168), .B2(n6146), .ZN(n6149)
         );
  NAND2_X1 U7124 ( .A1(n6167), .A2(REIP_REG_5__SCAN_IN), .ZN(n6148) );
  OAI211_X1 U7125 ( .C1(n6151), .C2(n6150), .A(n6149), .B(n6148), .ZN(U3013)
         );
  AOI21_X1 U7126 ( .B1(n6175), .B2(n6177), .A(n6172), .ZN(n6166) );
  INV_X1 U7127 ( .A(n6152), .ZN(n6153) );
  AOI222_X1 U7128 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6167), .B1(n6168), .B2(
        n6154), .C1(n6171), .C2(n6153), .ZN(n6158) );
  NOR2_X1 U7129 ( .A1(n6177), .A2(n6155), .ZN(n6162) );
  OAI211_X1 U7130 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6162), .B(n6156), .ZN(n6157) );
  OAI211_X1 U7131 ( .C1(n6166), .C2(n6159), .A(n6158), .B(n6157), .ZN(U3014)
         );
  AOI22_X1 U7132 ( .A1(n6168), .A2(n6160), .B1(n6167), .B2(REIP_REG_3__SCAN_IN), .ZN(n6164) );
  AOI22_X1 U7133 ( .A1(n6162), .A2(n6165), .B1(n6161), .B2(n6171), .ZN(n6163)
         );
  OAI211_X1 U7134 ( .C1(n6166), .C2(n6165), .A(n6164), .B(n6163), .ZN(U3015)
         );
  AOI22_X1 U7135 ( .A1(n6169), .A2(n6168), .B1(n6167), .B2(REIP_REG_2__SCAN_IN), .ZN(n6181) );
  AOI22_X1 U7136 ( .A1(n6172), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6171), 
        .B2(n6170), .ZN(n6180) );
  NAND3_X1 U7137 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6174), .A3(n6173), 
        .ZN(n6179) );
  OAI221_X1 U7138 ( .B1(n6177), .B2(n6176), .C1(n6177), .C2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(n6175), .ZN(n6178) );
  NAND4_X1 U7139 ( .A1(n6181), .A2(n6180), .A3(n6179), .A4(n6178), .ZN(U3016)
         );
  NOR2_X1 U7140 ( .A1(n6183), .A2(n6182), .ZN(U3019) );
  NAND3_X1 U7141 ( .A1(n6188), .A2(n6187), .A3(n6184), .ZN(n6251) );
  NOR2_X1 U7142 ( .A1(n6253), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6213)
         );
  AOI22_X1 U7143 ( .A1(n6304), .A2(n6213), .B1(n6212), .B2(n6185), .ZN(n6197)
         );
  NAND3_X1 U7144 ( .A1(n6188), .A2(n6187), .A3(n6186), .ZN(n6189) );
  NAND2_X1 U7145 ( .A1(n6189), .A2(n6500), .ZN(n6195) );
  AOI21_X1 U7146 ( .B1(n6190), .B2(n6256), .A(n6213), .ZN(n6194) );
  INV_X1 U7147 ( .A(n6194), .ZN(n6192) );
  NAND2_X1 U7148 ( .A1(n6308), .A2(n6193), .ZN(n6191) );
  OAI211_X1 U7149 ( .C1(n6195), .C2(n6192), .A(n6259), .B(n6191), .ZN(n6215)
         );
  OAI22_X1 U7150 ( .A1(n6195), .A2(n6194), .B1(n6193), .B2(n6405), .ZN(n6214)
         );
  AOI22_X1 U7151 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6215), .B1(n6303), 
        .B2(n6214), .ZN(n6196) );
  OAI211_X1 U7152 ( .C1(n6198), .C2(n6251), .A(n6197), .B(n6196), .ZN(U3044)
         );
  AOI22_X1 U7153 ( .A1(n6320), .A2(n6213), .B1(n6212), .B2(n6266), .ZN(n6200)
         );
  AOI22_X1 U7154 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6215), .B1(n6319), 
        .B2(n6214), .ZN(n6199) );
  OAI211_X1 U7155 ( .C1(n6269), .C2(n6251), .A(n6200), .B(n6199), .ZN(U3045)
         );
  AOI22_X1 U7156 ( .A1(n6326), .A2(n6213), .B1(n6212), .B2(n6270), .ZN(n6202)
         );
  AOI22_X1 U7157 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6215), .B1(n6325), 
        .B2(n6214), .ZN(n6201) );
  OAI211_X1 U7158 ( .C1(n6273), .C2(n6251), .A(n6202), .B(n6201), .ZN(U3046)
         );
  AOI22_X1 U7159 ( .A1(n6332), .A2(n6213), .B1(n6212), .B2(n6274), .ZN(n6204)
         );
  AOI22_X1 U7160 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6215), .B1(n6331), 
        .B2(n6214), .ZN(n6203) );
  OAI211_X1 U7161 ( .C1(n6277), .C2(n6251), .A(n6204), .B(n6203), .ZN(U3047)
         );
  AOI22_X1 U7162 ( .A1(n6338), .A2(n6213), .B1(n6212), .B2(n6278), .ZN(n6206)
         );
  AOI22_X1 U7163 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6215), .B1(n6337), 
        .B2(n6214), .ZN(n6205) );
  OAI211_X1 U7164 ( .C1(n6281), .C2(n6251), .A(n6206), .B(n6205), .ZN(U3048)
         );
  AOI22_X1 U7165 ( .A1(n6344), .A2(n6213), .B1(n6212), .B2(n6282), .ZN(n6208)
         );
  AOI22_X1 U7166 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6215), .B1(n6343), 
        .B2(n6214), .ZN(n6207) );
  OAI211_X1 U7167 ( .C1(n6285), .C2(n6251), .A(n6208), .B(n6207), .ZN(U3049)
         );
  AOI22_X1 U7168 ( .A1(n6350), .A2(n6213), .B1(n6212), .B2(n6286), .ZN(n6210)
         );
  AOI22_X1 U7169 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6215), .B1(n6349), 
        .B2(n6214), .ZN(n6209) );
  OAI211_X1 U7170 ( .C1(n6290), .C2(n6251), .A(n6210), .B(n6209), .ZN(U3050)
         );
  AOI22_X1 U7171 ( .A1(n6358), .A2(n6213), .B1(n6212), .B2(n6211), .ZN(n6217)
         );
  AOI22_X1 U7172 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6215), .B1(n6356), 
        .B2(n6214), .ZN(n6216) );
  OAI211_X1 U7173 ( .C1(n6218), .C2(n6251), .A(n6217), .B(n6216), .ZN(U3051)
         );
  NOR2_X1 U7174 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6219), .ZN(n6246)
         );
  NAND2_X1 U7175 ( .A1(n6310), .A2(n6500), .ZN(n6302) );
  INV_X1 U7176 ( .A(n6220), .ZN(n6221) );
  OAI22_X1 U7177 ( .A1(n6302), .A2(n6222), .B1(n6221), .B2(n6300), .ZN(n6245)
         );
  AOI22_X1 U7178 ( .A1(n6304), .A2(n6246), .B1(n6303), .B2(n6245), .ZN(n6232)
         );
  OAI22_X1 U7179 ( .A1(n6251), .A2(n6224), .B1(n6309), .B2(n6223), .ZN(n6229)
         );
  INV_X1 U7180 ( .A(n6246), .ZN(n6227) );
  AOI211_X1 U7181 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6227), .A(n6226), .B(
        n6225), .ZN(n6228) );
  OAI21_X1 U7182 ( .B1(n6230), .B2(n6229), .A(n6228), .ZN(n6248) );
  AOI22_X1 U7183 ( .A1(n6248), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n6315), 
        .B2(n6247), .ZN(n6231) );
  OAI211_X1 U7184 ( .C1(n6318), .C2(n6251), .A(n6232), .B(n6231), .ZN(U3052)
         );
  AOI22_X1 U7185 ( .A1(n6320), .A2(n6246), .B1(n6319), .B2(n6245), .ZN(n6234)
         );
  AOI22_X1 U7186 ( .A1(n6248), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n6321), 
        .B2(n6247), .ZN(n6233) );
  OAI211_X1 U7187 ( .C1(n6324), .C2(n6251), .A(n6234), .B(n6233), .ZN(U3053)
         );
  AOI22_X1 U7188 ( .A1(n6326), .A2(n6246), .B1(n6325), .B2(n6245), .ZN(n6236)
         );
  AOI22_X1 U7189 ( .A1(n6248), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n6327), 
        .B2(n6247), .ZN(n6235) );
  OAI211_X1 U7190 ( .C1(n6330), .C2(n6251), .A(n6236), .B(n6235), .ZN(U3054)
         );
  AOI22_X1 U7191 ( .A1(n6332), .A2(n6246), .B1(n6331), .B2(n6245), .ZN(n6238)
         );
  AOI22_X1 U7192 ( .A1(n6248), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6333), 
        .B2(n6247), .ZN(n6237) );
  OAI211_X1 U7193 ( .C1(n6336), .C2(n6251), .A(n6238), .B(n6237), .ZN(U3055)
         );
  AOI22_X1 U7194 ( .A1(n6338), .A2(n6246), .B1(n6337), .B2(n6245), .ZN(n6240)
         );
  AOI22_X1 U7195 ( .A1(n6248), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6339), 
        .B2(n6247), .ZN(n6239) );
  OAI211_X1 U7196 ( .C1(n6342), .C2(n6251), .A(n6240), .B(n6239), .ZN(U3056)
         );
  AOI22_X1 U7197 ( .A1(n6344), .A2(n6246), .B1(n6343), .B2(n6245), .ZN(n6242)
         );
  AOI22_X1 U7198 ( .A1(n6248), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n6345), 
        .B2(n6247), .ZN(n6241) );
  OAI211_X1 U7199 ( .C1(n6348), .C2(n6251), .A(n6242), .B(n6241), .ZN(U3057)
         );
  AOI22_X1 U7200 ( .A1(n6350), .A2(n6246), .B1(n6349), .B2(n6245), .ZN(n6244)
         );
  AOI22_X1 U7201 ( .A1(n6248), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6351), 
        .B2(n6247), .ZN(n6243) );
  OAI211_X1 U7202 ( .C1(n6354), .C2(n6251), .A(n6244), .B(n6243), .ZN(U3058)
         );
  AOI22_X1 U7203 ( .A1(n6358), .A2(n6246), .B1(n6356), .B2(n6245), .ZN(n6250)
         );
  AOI22_X1 U7204 ( .A1(n6248), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n6360), 
        .B2(n6247), .ZN(n6249) );
  OAI211_X1 U7205 ( .C1(n6365), .C2(n6251), .A(n6250), .B(n6249), .ZN(U3059)
         );
  INV_X1 U7206 ( .A(n6364), .ZN(n6292) );
  NOR2_X1 U7207 ( .A1(n6253), .A2(n6383), .ZN(n6291) );
  AOI22_X1 U7208 ( .A1(n6315), .A2(n6292), .B1(n6304), .B2(n6291), .ZN(n6265)
         );
  OAI21_X1 U7209 ( .B1(n6255), .B2(n6254), .A(n6500), .ZN(n6263) );
  AOI21_X1 U7210 ( .B1(n6257), .B2(n6256), .A(n6291), .ZN(n6262) );
  INV_X1 U7211 ( .A(n6262), .ZN(n6260) );
  NAND2_X1 U7212 ( .A1(n6308), .A2(n6261), .ZN(n6258) );
  OAI211_X1 U7213 ( .C1(n6263), .C2(n6260), .A(n6259), .B(n6258), .ZN(n6294)
         );
  OAI22_X1 U7214 ( .A1(n6263), .A2(n6262), .B1(n6261), .B2(n6405), .ZN(n6293)
         );
  AOI22_X1 U7215 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6294), .B1(n6303), 
        .B2(n6293), .ZN(n6264) );
  OAI211_X1 U7216 ( .C1(n6318), .C2(n6297), .A(n6265), .B(n6264), .ZN(U3108)
         );
  INV_X1 U7217 ( .A(n6297), .ZN(n6287) );
  AOI22_X1 U7218 ( .A1(n6287), .A2(n6266), .B1(n6320), .B2(n6291), .ZN(n6268)
         );
  AOI22_X1 U7219 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6294), .B1(n6319), 
        .B2(n6293), .ZN(n6267) );
  OAI211_X1 U7220 ( .C1(n6269), .C2(n6364), .A(n6268), .B(n6267), .ZN(U3109)
         );
  AOI22_X1 U7221 ( .A1(n6287), .A2(n6270), .B1(n6326), .B2(n6291), .ZN(n6272)
         );
  AOI22_X1 U7222 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6294), .B1(n6325), 
        .B2(n6293), .ZN(n6271) );
  OAI211_X1 U7223 ( .C1(n6273), .C2(n6364), .A(n6272), .B(n6271), .ZN(U3110)
         );
  AOI22_X1 U7224 ( .A1(n6287), .A2(n6274), .B1(n6332), .B2(n6291), .ZN(n6276)
         );
  AOI22_X1 U7225 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6294), .B1(n6331), 
        .B2(n6293), .ZN(n6275) );
  OAI211_X1 U7226 ( .C1(n6277), .C2(n6364), .A(n6276), .B(n6275), .ZN(U3111)
         );
  AOI22_X1 U7227 ( .A1(n6287), .A2(n6278), .B1(n6338), .B2(n6291), .ZN(n6280)
         );
  AOI22_X1 U7228 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6294), .B1(n6337), 
        .B2(n6293), .ZN(n6279) );
  OAI211_X1 U7229 ( .C1(n6281), .C2(n6364), .A(n6280), .B(n6279), .ZN(U3112)
         );
  AOI22_X1 U7230 ( .A1(n6287), .A2(n6282), .B1(n6344), .B2(n6291), .ZN(n6284)
         );
  AOI22_X1 U7231 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6294), .B1(n6343), 
        .B2(n6293), .ZN(n6283) );
  OAI211_X1 U7232 ( .C1(n6285), .C2(n6364), .A(n6284), .B(n6283), .ZN(U3113)
         );
  AOI22_X1 U7233 ( .A1(n6287), .A2(n6286), .B1(n6350), .B2(n6291), .ZN(n6289)
         );
  AOI22_X1 U7234 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6294), .B1(n6349), 
        .B2(n6293), .ZN(n6288) );
  OAI211_X1 U7235 ( .C1(n6290), .C2(n6364), .A(n6289), .B(n6288), .ZN(U3114)
         );
  AOI22_X1 U7236 ( .A1(n6360), .A2(n6292), .B1(n6358), .B2(n6291), .ZN(n6296)
         );
  AOI22_X1 U7237 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6294), .B1(n6356), 
        .B2(n6293), .ZN(n6295) );
  OAI211_X1 U7238 ( .C1(n6365), .C2(n6297), .A(n6296), .B(n6295), .ZN(U3115)
         );
  NOR2_X1 U7239 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6298), .ZN(n6357)
         );
  OAI22_X1 U7240 ( .A1(n6302), .A2(n6301), .B1(n6300), .B2(n6299), .ZN(n6355)
         );
  AOI22_X1 U7241 ( .A1(n6304), .A2(n6357), .B1(n6303), .B2(n6355), .ZN(n6317)
         );
  INV_X1 U7242 ( .A(n6359), .ZN(n6306) );
  AOI21_X1 U7243 ( .B1(n6306), .B2(n6364), .A(n6305), .ZN(n6307) );
  AOI211_X1 U7244 ( .C1(n6310), .C2(n6309), .A(n6308), .B(n6307), .ZN(n6314)
         );
  OAI211_X1 U7245 ( .C1(n6483), .C2(n6357), .A(n6312), .B(n6311), .ZN(n6313)
         );
  AOI22_X1 U7246 ( .A1(n6361), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n6315), 
        .B2(n6359), .ZN(n6316) );
  OAI211_X1 U7247 ( .C1(n6318), .C2(n6364), .A(n6317), .B(n6316), .ZN(U3116)
         );
  AOI22_X1 U7248 ( .A1(n6320), .A2(n6357), .B1(n6319), .B2(n6355), .ZN(n6323)
         );
  AOI22_X1 U7249 ( .A1(n6361), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n6321), 
        .B2(n6359), .ZN(n6322) );
  OAI211_X1 U7250 ( .C1(n6324), .C2(n6364), .A(n6323), .B(n6322), .ZN(U3117)
         );
  AOI22_X1 U7251 ( .A1(n6326), .A2(n6357), .B1(n6325), .B2(n6355), .ZN(n6329)
         );
  AOI22_X1 U7252 ( .A1(n6361), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n6327), 
        .B2(n6359), .ZN(n6328) );
  OAI211_X1 U7253 ( .C1(n6330), .C2(n6364), .A(n6329), .B(n6328), .ZN(U3118)
         );
  AOI22_X1 U7254 ( .A1(n6332), .A2(n6357), .B1(n6331), .B2(n6355), .ZN(n6335)
         );
  AOI22_X1 U7255 ( .A1(n6361), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n6333), 
        .B2(n6359), .ZN(n6334) );
  OAI211_X1 U7256 ( .C1(n6336), .C2(n6364), .A(n6335), .B(n6334), .ZN(U3119)
         );
  AOI22_X1 U7257 ( .A1(n6338), .A2(n6357), .B1(n6337), .B2(n6355), .ZN(n6341)
         );
  AOI22_X1 U7258 ( .A1(n6361), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n6339), 
        .B2(n6359), .ZN(n6340) );
  OAI211_X1 U7259 ( .C1(n6342), .C2(n6364), .A(n6341), .B(n6340), .ZN(U3120)
         );
  AOI22_X1 U7260 ( .A1(n6344), .A2(n6357), .B1(n6343), .B2(n6355), .ZN(n6347)
         );
  AOI22_X1 U7261 ( .A1(n6361), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n6345), 
        .B2(n6359), .ZN(n6346) );
  OAI211_X1 U7262 ( .C1(n6348), .C2(n6364), .A(n6347), .B(n6346), .ZN(U3121)
         );
  AOI22_X1 U7263 ( .A1(n6350), .A2(n6357), .B1(n6349), .B2(n6355), .ZN(n6353)
         );
  AOI22_X1 U7264 ( .A1(n6361), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6351), 
        .B2(n6359), .ZN(n6352) );
  OAI211_X1 U7265 ( .C1(n6354), .C2(n6364), .A(n6353), .B(n6352), .ZN(U3122)
         );
  AOI22_X1 U7266 ( .A1(n6358), .A2(n6357), .B1(n6356), .B2(n6355), .ZN(n6363)
         );
  AOI22_X1 U7267 ( .A1(n6361), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6360), 
        .B2(n6359), .ZN(n6362) );
  OAI211_X1 U7268 ( .C1(n6365), .C2(n6364), .A(n6363), .B(n6362), .ZN(U3123)
         );
  INV_X1 U7269 ( .A(n6385), .ZN(n6382) );
  INV_X1 U7270 ( .A(n6366), .ZN(n6368) );
  OAI211_X1 U7271 ( .C1(n6369), .C2(n6368), .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n6367), .ZN(n6371) );
  OAI21_X1 U7272 ( .B1(n6372), .B2(n6371), .A(n6370), .ZN(n6374) );
  NAND2_X1 U7273 ( .A1(n6372), .A2(n6371), .ZN(n6373) );
  OAI21_X1 U7274 ( .B1(n6375), .B2(n6374), .A(n6373), .ZN(n6377) );
  NAND2_X1 U7275 ( .A1(n6376), .A2(n6377), .ZN(n6379) );
  INV_X1 U7276 ( .A(n6377), .ZN(n6378) );
  AOI22_X1 U7277 ( .A1(n6380), .A2(n6379), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6378), .ZN(n6381) );
  AOI21_X1 U7278 ( .B1(n6383), .B2(n6382), .A(n6381), .ZN(n6384) );
  AOI211_X1 U7279 ( .C1(n6385), .C2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n6384), .ZN(n6394) );
  INV_X1 U7280 ( .A(n6386), .ZN(n6393) );
  NOR2_X1 U7281 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6390) );
  OAI211_X1 U7282 ( .C1(n6390), .C2(n6389), .A(n6388), .B(n6387), .ZN(n6391)
         );
  NOR4_X1 U7283 ( .A1(n6394), .A2(n6393), .A3(n6392), .A4(n6391), .ZN(n6404)
         );
  INV_X1 U7284 ( .A(n6404), .ZN(n6396) );
  OAI22_X1 U7285 ( .A1(n6396), .A2(n6407), .B1(n6592), .B2(n6395), .ZN(n6397)
         );
  OAI21_X1 U7286 ( .B1(n6399), .B2(n6398), .A(n6397), .ZN(n6482) );
  OAI21_X1 U7287 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6592), .A(n6482), .ZN(
        n6406) );
  AOI221_X1 U7288 ( .B1(n6401), .B2(STATE2_REG_0__SCAN_IN), .C1(n6406), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6400), .ZN(n6403) );
  OAI211_X1 U7289 ( .C1(n6413), .C2(n6484), .A(n6520), .B(n6482), .ZN(n6402)
         );
  OAI211_X1 U7290 ( .C1(n6404), .C2(n6407), .A(n6403), .B(n6402), .ZN(U3148)
         );
  NAND2_X1 U7291 ( .A1(n6520), .A2(n6405), .ZN(n6414) );
  NAND3_X1 U7292 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6414), .A3(n6406), .ZN(
        n6412) );
  OAI21_X1 U7293 ( .B1(READY_N), .B2(n6408), .A(n6407), .ZN(n6410) );
  AOI21_X1 U7294 ( .B1(n6410), .B2(n6482), .A(n6409), .ZN(n6411) );
  NAND2_X1 U7295 ( .A1(n6412), .A2(n6411), .ZN(U3149) );
  INV_X1 U7296 ( .A(n6413), .ZN(n6507) );
  OAI211_X1 U7297 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6592), .A(n6480), .B(
        n6414), .ZN(n6416) );
  OAI21_X1 U7298 ( .B1(n6507), .B2(n6416), .A(n6415), .ZN(U3150) );
  INV_X1 U7299 ( .A(n6479), .ZN(n6475) );
  AND2_X1 U7300 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6475), .ZN(U3151) );
  AND2_X1 U7301 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6475), .ZN(U3152) );
  AND2_X1 U7302 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6475), .ZN(U3153) );
  AND2_X1 U7303 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6475), .ZN(U3154) );
  INV_X1 U7304 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6595) );
  NOR2_X1 U7305 ( .A1(n6479), .A2(n6595), .ZN(U3155) );
  INV_X1 U7306 ( .A(DATAWIDTH_REG_26__SCAN_IN), .ZN(n6628) );
  NOR2_X1 U7307 ( .A1(n6479), .A2(n6628), .ZN(U3156) );
  AND2_X1 U7308 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6475), .ZN(U3157) );
  AND2_X1 U7309 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6475), .ZN(U3158) );
  AND2_X1 U7310 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6475), .ZN(U3159) );
  AND2_X1 U7311 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6475), .ZN(U3160) );
  INV_X1 U7312 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6518) );
  NOR2_X1 U7313 ( .A1(n6479), .A2(n6518), .ZN(U3161) );
  AND2_X1 U7314 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6475), .ZN(U3162) );
  AND2_X1 U7315 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6475), .ZN(U3163) );
  AND2_X1 U7316 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6475), .ZN(U3164) );
  AND2_X1 U7317 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6475), .ZN(U3165) );
  INV_X1 U7318 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6536) );
  NOR2_X1 U7319 ( .A1(n6479), .A2(n6536), .ZN(U3166) );
  AND2_X1 U7320 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6475), .ZN(U3167) );
  AND2_X1 U7321 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6475), .ZN(U3168) );
  AND2_X1 U7322 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6475), .ZN(U3169) );
  AND2_X1 U7323 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6475), .ZN(U3170) );
  AND2_X1 U7324 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6475), .ZN(U3171) );
  AND2_X1 U7325 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6475), .ZN(U3172) );
  AND2_X1 U7326 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6475), .ZN(U3173) );
  AND2_X1 U7327 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6475), .ZN(U3174) );
  AND2_X1 U7328 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6475), .ZN(U3175) );
  AND2_X1 U7329 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6475), .ZN(U3176) );
  AND2_X1 U7330 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6475), .ZN(U3177) );
  INV_X1 U7331 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6612) );
  NOR2_X1 U7332 ( .A1(n6479), .A2(n6612), .ZN(U3178) );
  AND2_X1 U7333 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6475), .ZN(U3179) );
  AND2_X1 U7334 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6475), .ZN(U3180) );
  INV_X1 U7335 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6423) );
  NOR2_X1 U7336 ( .A1(n6548), .A2(n6423), .ZN(n6426) );
  AOI22_X1 U7337 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6430) );
  AND2_X1 U7338 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6420) );
  INV_X2 U7339 ( .A(n6512), .ZN(n6663) );
  INV_X1 U7340 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6418) );
  INV_X1 U7341 ( .A(NA_N), .ZN(n6427) );
  AOI211_X1 U7342 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6427), .A(
        STATE_REG_0__SCAN_IN), .B(n6426), .ZN(n6432) );
  AOI221_X1 U7343 ( .B1(n6420), .B2(n6663), .C1(n6418), .C2(n6663), .A(n6432), 
        .ZN(n6417) );
  OAI21_X1 U7344 ( .B1(n6426), .B2(n6430), .A(n6417), .ZN(U3181) );
  NOR2_X1 U7345 ( .A1(n6424), .A2(n6418), .ZN(n6428) );
  NAND2_X1 U7346 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6419) );
  OAI21_X1 U7347 ( .B1(n6428), .B2(n6420), .A(n6419), .ZN(n6421) );
  OAI211_X1 U7348 ( .C1(n6423), .C2(n6592), .A(n6422), .B(n6421), .ZN(U3182)
         );
  AOI221_X1 U7349 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6592), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6425) );
  AOI221_X1 U7350 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6425), .C2(HOLD), .A(n6424), .ZN(n6431) );
  AOI21_X1 U7351 ( .B1(n6428), .B2(n6427), .A(n6426), .ZN(n6429) );
  OAI22_X1 U7352 ( .A1(n6432), .A2(n6431), .B1(n6430), .B2(n6429), .ZN(U3183)
         );
  NOR2_X2 U7353 ( .A1(n6548), .A2(n6663), .ZN(n6662) );
  INV_X1 U7354 ( .A(n6662), .ZN(n6472) );
  NOR2_X2 U7355 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6663), .ZN(n6661) );
  AOI22_X1 U7356 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6661), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6663), .ZN(n6433) );
  OAI21_X1 U7357 ( .B1(n6490), .B2(n6472), .A(n6433), .ZN(U3184) );
  INV_X1 U7358 ( .A(n6661), .ZN(n6466) );
  AOI22_X1 U7359 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6662), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6663), .ZN(n6434) );
  OAI21_X1 U7360 ( .B1(n6529), .B2(n6466), .A(n6434), .ZN(U3185) );
  AOI22_X1 U7361 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6662), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6663), .ZN(n6435) );
  OAI21_X1 U7362 ( .B1(n6436), .B2(n6466), .A(n6435), .ZN(U3186) );
  AOI22_X1 U7363 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6662), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6663), .ZN(n6437) );
  OAI21_X1 U7364 ( .B1(n4459), .B2(n6466), .A(n6437), .ZN(U3187) );
  AOI22_X1 U7365 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6661), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6663), .ZN(n6438) );
  OAI21_X1 U7366 ( .B1(n4459), .B2(n6472), .A(n6438), .ZN(U3188) );
  AOI22_X1 U7367 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6661), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6663), .ZN(n6439) );
  OAI21_X1 U7368 ( .B1(n6554), .B2(n6472), .A(n6439), .ZN(U3190) );
  AOI22_X1 U7369 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6662), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6663), .ZN(n6440) );
  OAI21_X1 U7370 ( .B1(n4907), .B2(n6466), .A(n6440), .ZN(U3191) );
  INV_X1 U7371 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6545) );
  OAI222_X1 U7372 ( .A1(n6472), .A2(n4907), .B1(n6545), .B2(n6512), .C1(n6442), 
        .C2(n6466), .ZN(U3192) );
  AOI22_X1 U7373 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6661), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6663), .ZN(n6441) );
  OAI21_X1 U7374 ( .B1(n6442), .B2(n6472), .A(n6441), .ZN(U3193) );
  AOI22_X1 U7375 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6662), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6663), .ZN(n6443) );
  OAI21_X1 U7376 ( .B1(n6445), .B2(n6466), .A(n6443), .ZN(U3194) );
  AOI22_X1 U7377 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6661), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6663), .ZN(n6444) );
  OAI21_X1 U7378 ( .B1(n6445), .B2(n6472), .A(n6444), .ZN(U3195) );
  AOI22_X1 U7379 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6662), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6663), .ZN(n6446) );
  OAI21_X1 U7380 ( .B1(n6448), .B2(n6466), .A(n6446), .ZN(U3196) );
  AOI22_X1 U7381 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6661), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6663), .ZN(n6447) );
  OAI21_X1 U7382 ( .B1(n6448), .B2(n6472), .A(n6447), .ZN(U3197) );
  AOI22_X1 U7383 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6662), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6663), .ZN(n6449) );
  OAI21_X1 U7384 ( .B1(n6451), .B2(n6466), .A(n6449), .ZN(U3198) );
  AOI22_X1 U7385 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6661), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6663), .ZN(n6450) );
  OAI21_X1 U7386 ( .B1(n6451), .B2(n6472), .A(n6450), .ZN(U3199) );
  AOI22_X1 U7387 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6662), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6663), .ZN(n6452) );
  OAI21_X1 U7388 ( .B1(n6453), .B2(n6466), .A(n6452), .ZN(U3200) );
  AOI22_X1 U7389 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6662), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6663), .ZN(n6454) );
  OAI21_X1 U7390 ( .B1(n5084), .B2(n6466), .A(n6454), .ZN(U3201) );
  AOI22_X1 U7391 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6661), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6663), .ZN(n6455) );
  OAI21_X1 U7392 ( .B1(n5084), .B2(n6472), .A(n6455), .ZN(U3202) );
  INV_X1 U7393 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6530) );
  OAI222_X1 U7394 ( .A1(n6472), .A2(n5110), .B1(n6530), .B2(n6512), .C1(n6457), 
        .C2(n6466), .ZN(U3203) );
  AOI22_X1 U7395 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6661), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6663), .ZN(n6456) );
  OAI21_X1 U7396 ( .B1(n6457), .B2(n6472), .A(n6456), .ZN(U3204) );
  AOI22_X1 U7397 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6662), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6663), .ZN(n6458) );
  OAI21_X1 U7398 ( .B1(n5259), .B2(n6466), .A(n6458), .ZN(U3205) );
  AOI22_X1 U7399 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6661), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6663), .ZN(n6459) );
  OAI21_X1 U7400 ( .B1(n5259), .B2(n6472), .A(n6459), .ZN(U3206) );
  AOI22_X1 U7401 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6662), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6663), .ZN(n6460) );
  OAI21_X1 U7402 ( .B1(n6462), .B2(n6466), .A(n6460), .ZN(U3207) );
  AOI22_X1 U7403 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6661), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6663), .ZN(n6461) );
  OAI21_X1 U7404 ( .B1(n6462), .B2(n6472), .A(n6461), .ZN(U3208) );
  AOI22_X1 U7405 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6662), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6663), .ZN(n6463) );
  OAI21_X1 U7406 ( .B1(n6464), .B2(n6466), .A(n6463), .ZN(U3209) );
  AOI22_X1 U7407 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6662), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6663), .ZN(n6465) );
  OAI21_X1 U7408 ( .B1(n6468), .B2(n6466), .A(n6465), .ZN(U3210) );
  AOI22_X1 U7409 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6661), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6663), .ZN(n6467) );
  OAI21_X1 U7410 ( .B1(n6468), .B2(n6472), .A(n6467), .ZN(U3211) );
  AOI22_X1 U7411 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6661), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6663), .ZN(n6469) );
  OAI21_X1 U7412 ( .B1(n6470), .B2(n6472), .A(n6469), .ZN(U3212) );
  AOI22_X1 U7413 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6661), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6663), .ZN(n6471) );
  OAI21_X1 U7414 ( .B1(n6473), .B2(n6472), .A(n6471), .ZN(U3213) );
  MUX2_X1 U7415 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6512), .Z(U3445) );
  MUX2_X1 U7416 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6512), .Z(U3446) );
  MUX2_X1 U7417 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6512), .Z(U3447) );
  MUX2_X1 U7418 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6512), .Z(U3448) );
  INV_X1 U7419 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6476) );
  INV_X1 U7420 ( .A(n6477), .ZN(n6474) );
  AOI21_X1 U7421 ( .B1(n6476), .B2(n6475), .A(n6474), .ZN(U3451) );
  OAI21_X1 U7422 ( .B1(n6479), .B2(n6478), .A(n6477), .ZN(U3452) );
  OAI211_X1 U7423 ( .C1(n6483), .C2(n6482), .A(n6481), .B(n6480), .ZN(U3453)
         );
  OAI22_X1 U7424 ( .A1(n6487), .A2(n6486), .B1(n6485), .B2(n6484), .ZN(n6489)
         );
  MUX2_X1 U7425 ( .A(n6489), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6488), 
        .Z(U3456) );
  AOI21_X1 U7426 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6491) );
  AOI22_X1 U7427 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6491), .B2(n6490), .ZN(n6494) );
  INV_X1 U7428 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6493) );
  AOI22_X1 U7429 ( .A1(n6497), .A2(n6494), .B1(n6493), .B2(n6492), .ZN(U3468)
         );
  INV_X1 U7430 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6496) );
  OAI21_X1 U7431 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6497), .ZN(n6495) );
  OAI21_X1 U7432 ( .B1(n6497), .B2(n6496), .A(n6495), .ZN(U3469) );
  NAND2_X1 U7433 ( .A1(n6663), .A2(W_R_N_REG_SCAN_IN), .ZN(n6498) );
  OAI21_X1 U7434 ( .B1(n6663), .B2(READREQUEST_REG_SCAN_IN), .A(n6498), .ZN(
        U3470) );
  AOI211_X1 U7435 ( .C1(n6592), .C2(n6501), .A(n6500), .B(n6499), .ZN(n6502)
         );
  AND2_X1 U7436 ( .A1(n6503), .A2(n6502), .ZN(n6511) );
  INV_X1 U7437 ( .A(n6504), .ZN(n6505) );
  OAI211_X1 U7438 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6506), .A(n6505), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6508) );
  AOI21_X1 U7439 ( .B1(n6508), .B2(STATE2_REG_0__SCAN_IN), .A(n6507), .ZN(
        n6510) );
  NAND2_X1 U7440 ( .A1(n6511), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6509) );
  OAI21_X1 U7441 ( .B1(n6511), .B2(n6510), .A(n6509), .ZN(U3472) );
  MUX2_X1 U7442 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6512), .Z(U3473) );
  INV_X1 U7443 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n6514) );
  AOI22_X1 U7444 ( .A1(n6515), .A2(keyinput28), .B1(n6514), .B2(keyinput63), 
        .ZN(n6513) );
  OAI221_X1 U7445 ( .B1(n6515), .B2(keyinput28), .C1(n6514), .C2(keyinput63), 
        .A(n6513), .ZN(n6527) );
  INV_X1 U7446 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n6517) );
  AOI22_X1 U7447 ( .A1(n6518), .A2(keyinput49), .B1(n6517), .B2(keyinput24), 
        .ZN(n6516) );
  OAI221_X1 U7448 ( .B1(n6518), .B2(keyinput49), .C1(n6517), .C2(keyinput24), 
        .A(n6516), .ZN(n6526) );
  AOI22_X1 U7449 ( .A1(n3007), .A2(keyinput56), .B1(n6520), .B2(keyinput4), 
        .ZN(n6519) );
  OAI221_X1 U7450 ( .B1(n3007), .B2(keyinput56), .C1(n6520), .C2(keyinput4), 
        .A(n6519), .ZN(n6525) );
  INV_X1 U7451 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n6523) );
  INV_X1 U7452 ( .A(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n6522) );
  AOI22_X1 U7453 ( .A1(n6523), .A2(keyinput60), .B1(n6522), .B2(keyinput2), 
        .ZN(n6521) );
  OAI221_X1 U7454 ( .B1(n6523), .B2(keyinput60), .C1(n6522), .C2(keyinput2), 
        .A(n6521), .ZN(n6524) );
  NOR4_X1 U7455 ( .A1(n6527), .A2(n6526), .A3(n6525), .A4(n6524), .ZN(n6577)
         );
  AOI22_X1 U7456 ( .A1(n6530), .A2(keyinput47), .B1(n6529), .B2(keyinput41), 
        .ZN(n6528) );
  OAI221_X1 U7457 ( .B1(n6530), .B2(keyinput47), .C1(n6529), .C2(keyinput41), 
        .A(n6528), .ZN(n6543) );
  AOI22_X1 U7458 ( .A1(n6533), .A2(keyinput7), .B1(keyinput57), .B2(n6532), 
        .ZN(n6531) );
  OAI221_X1 U7459 ( .B1(n6533), .B2(keyinput7), .C1(n6532), .C2(keyinput57), 
        .A(n6531), .ZN(n6542) );
  INV_X1 U7460 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6535) );
  AOI22_X1 U7461 ( .A1(n6536), .A2(keyinput20), .B1(n6535), .B2(keyinput53), 
        .ZN(n6534) );
  OAI221_X1 U7462 ( .B1(n6536), .B2(keyinput20), .C1(n6535), .C2(keyinput53), 
        .A(n6534), .ZN(n6541) );
  XOR2_X1 U7463 ( .A(n6537), .B(keyinput15), .Z(n6539) );
  XNOR2_X1 U7464 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .B(keyinput37), .ZN(n6538)
         );
  NAND2_X1 U7465 ( .A1(n6539), .A2(n6538), .ZN(n6540) );
  NOR4_X1 U7466 ( .A1(n6543), .A2(n6542), .A3(n6541), .A4(n6540), .ZN(n6576)
         );
  INV_X1 U7467 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n6546) );
  AOI22_X1 U7468 ( .A1(n6546), .A2(keyinput32), .B1(keyinput38), .B2(n6545), 
        .ZN(n6544) );
  OAI221_X1 U7469 ( .B1(n6546), .B2(keyinput32), .C1(n6545), .C2(keyinput38), 
        .A(n6544), .ZN(n6559) );
  AOI22_X1 U7470 ( .A1(n6549), .A2(keyinput22), .B1(n6548), .B2(keyinput51), 
        .ZN(n6547) );
  OAI221_X1 U7471 ( .B1(n6549), .B2(keyinput22), .C1(n6548), .C2(keyinput51), 
        .A(n6547), .ZN(n6558) );
  AOI22_X1 U7472 ( .A1(n6552), .A2(keyinput34), .B1(n6551), .B2(keyinput35), 
        .ZN(n6550) );
  OAI221_X1 U7473 ( .B1(n6552), .B2(keyinput34), .C1(n6551), .C2(keyinput35), 
        .A(n6550), .ZN(n6557) );
  INV_X1 U7474 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n6555) );
  AOI22_X1 U7475 ( .A1(n6555), .A2(keyinput55), .B1(n6554), .B2(keyinput8), 
        .ZN(n6553) );
  OAI221_X1 U7476 ( .B1(n6555), .B2(keyinput55), .C1(n6554), .C2(keyinput8), 
        .A(n6553), .ZN(n6556) );
  NOR4_X1 U7477 ( .A1(n6559), .A2(n6558), .A3(n6557), .A4(n6556), .ZN(n6575)
         );
  AOI22_X1 U7478 ( .A1(n3765), .A2(keyinput52), .B1(keyinput39), .B2(n6561), 
        .ZN(n6560) );
  OAI221_X1 U7479 ( .B1(n3765), .B2(keyinput52), .C1(n6561), .C2(keyinput39), 
        .A(n6560), .ZN(n6573) );
  INV_X1 U7480 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6564) );
  INV_X1 U7481 ( .A(DATAI_30_), .ZN(n6563) );
  AOI22_X1 U7482 ( .A1(n6564), .A2(keyinput26), .B1(keyinput33), .B2(n6563), 
        .ZN(n6562) );
  OAI221_X1 U7483 ( .B1(n6564), .B2(keyinput26), .C1(n6563), .C2(keyinput33), 
        .A(n6562), .ZN(n6572) );
  INV_X1 U7484 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6567) );
  OAI221_X1 U7485 ( .B1(n6567), .B2(keyinput48), .C1(n6566), .C2(keyinput18), 
        .A(n6565), .ZN(n6571) );
  XNOR2_X1 U7486 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .B(keyinput30), .ZN(n6569)
         );
  XNOR2_X1 U7487 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .B(keyinput23), .ZN(n6568) );
  NAND2_X1 U7488 ( .A1(n6569), .A2(n6568), .ZN(n6570) );
  NOR4_X1 U7489 ( .A1(n6573), .A2(n6572), .A3(n6571), .A4(n6570), .ZN(n6574)
         );
  NAND4_X1 U7490 ( .A1(n6577), .A2(n6576), .A3(n6575), .A4(n6574), .ZN(n6639)
         );
  AOI22_X1 U7491 ( .A1(n3904), .A2(keyinput43), .B1(n6579), .B2(keyinput16), 
        .ZN(n6578) );
  OAI221_X1 U7492 ( .B1(n3904), .B2(keyinput43), .C1(n6579), .C2(keyinput16), 
        .A(n6578), .ZN(n6590) );
  AOI22_X1 U7493 ( .A1(n6581), .A2(keyinput54), .B1(n4880), .B2(keyinput61), 
        .ZN(n6580) );
  OAI221_X1 U7494 ( .B1(n6581), .B2(keyinput54), .C1(n4880), .C2(keyinput61), 
        .A(n6580), .ZN(n6589) );
  AOI22_X1 U7495 ( .A1(n6584), .A2(keyinput58), .B1(keyinput44), .B2(n6583), 
        .ZN(n6582) );
  OAI221_X1 U7496 ( .B1(n6584), .B2(keyinput58), .C1(n6583), .C2(keyinput44), 
        .A(n6582), .ZN(n6588) );
  AOI22_X1 U7497 ( .A1(n3690), .A2(keyinput10), .B1(n6586), .B2(keyinput29), 
        .ZN(n6585) );
  OAI221_X1 U7498 ( .B1(n3690), .B2(keyinput10), .C1(n6586), .C2(keyinput29), 
        .A(n6585), .ZN(n6587) );
  NOR4_X1 U7499 ( .A1(n6590), .A2(n6589), .A3(n6588), .A4(n6587), .ZN(n6637)
         );
  AOI22_X1 U7500 ( .A1(n4309), .A2(keyinput46), .B1(n6592), .B2(keyinput9), 
        .ZN(n6591) );
  OAI221_X1 U7501 ( .B1(n4309), .B2(keyinput46), .C1(n6592), .C2(keyinput9), 
        .A(n6591), .ZN(n6604) );
  AOI22_X1 U7502 ( .A1(n6595), .A2(keyinput27), .B1(n6594), .B2(keyinput59), 
        .ZN(n6593) );
  OAI221_X1 U7503 ( .B1(n6595), .B2(keyinput27), .C1(n6594), .C2(keyinput59), 
        .A(n6593), .ZN(n6603) );
  AOI22_X1 U7504 ( .A1(n6597), .A2(keyinput0), .B1(n6057), .B2(keyinput5), 
        .ZN(n6596) );
  OAI221_X1 U7505 ( .B1(n6597), .B2(keyinput0), .C1(n6057), .C2(keyinput5), 
        .A(n6596), .ZN(n6602) );
  INV_X1 U7506 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n6598) );
  XOR2_X1 U7507 ( .A(n6598), .B(keyinput50), .Z(n6600) );
  XNOR2_X1 U7508 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(keyinput31), .ZN(
        n6599) );
  NAND2_X1 U7509 ( .A1(n6600), .A2(n6599), .ZN(n6601) );
  NOR4_X1 U7510 ( .A1(n6604), .A2(n6603), .A3(n6602), .A4(n6601), .ZN(n6636)
         );
  INV_X1 U7511 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n6606) );
  AOI22_X1 U7512 ( .A1(n6607), .A2(keyinput62), .B1(keyinput6), .B2(n6606), 
        .ZN(n6605) );
  OAI221_X1 U7513 ( .B1(n6607), .B2(keyinput62), .C1(n6606), .C2(keyinput6), 
        .A(n6605), .ZN(n6618) );
  AOI22_X1 U7514 ( .A1(n5787), .A2(keyinput21), .B1(keyinput13), .B2(n6609), 
        .ZN(n6608) );
  OAI221_X1 U7515 ( .B1(n5787), .B2(keyinput21), .C1(n6609), .C2(keyinput13), 
        .A(n6608), .ZN(n6617) );
  INV_X1 U7516 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n6611) );
  AOI22_X1 U7517 ( .A1(n6612), .A2(keyinput45), .B1(n6611), .B2(keyinput25), 
        .ZN(n6610) );
  OAI221_X1 U7518 ( .B1(n6612), .B2(keyinput45), .C1(n6611), .C2(keyinput25), 
        .A(n6610), .ZN(n6616) );
  AOI22_X1 U7519 ( .A1(n5579), .A2(keyinput17), .B1(keyinput1), .B2(n6614), 
        .ZN(n6613) );
  OAI221_X1 U7520 ( .B1(n5579), .B2(keyinput17), .C1(n6614), .C2(keyinput1), 
        .A(n6613), .ZN(n6615) );
  NOR4_X1 U7521 ( .A1(n6618), .A2(n6617), .A3(n6616), .A4(n6615), .ZN(n6635)
         );
  INV_X1 U7522 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n6621) );
  INV_X1 U7523 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6620) );
  AOI22_X1 U7524 ( .A1(n6621), .A2(keyinput14), .B1(n6620), .B2(keyinput12), 
        .ZN(n6619) );
  OAI221_X1 U7525 ( .B1(n6621), .B2(keyinput14), .C1(n6620), .C2(keyinput12), 
        .A(n6619), .ZN(n6633) );
  AOI22_X1 U7526 ( .A1(n3036), .A2(keyinput40), .B1(keyinput11), .B2(n6623), 
        .ZN(n6622) );
  OAI221_X1 U7527 ( .B1(n3036), .B2(keyinput40), .C1(n6623), .C2(keyinput11), 
        .A(n6622), .ZN(n6632) );
  INV_X1 U7528 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n6626) );
  AOI22_X1 U7529 ( .A1(n6626), .A2(keyinput3), .B1(keyinput42), .B2(n6625), 
        .ZN(n6624) );
  OAI221_X1 U7530 ( .B1(n6626), .B2(keyinput3), .C1(n6625), .C2(keyinput42), 
        .A(n6624), .ZN(n6631) );
  INV_X1 U7531 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n6629) );
  AOI22_X1 U7532 ( .A1(n6629), .A2(keyinput19), .B1(keyinput36), .B2(n6628), 
        .ZN(n6627) );
  OAI221_X1 U7533 ( .B1(n6629), .B2(keyinput19), .C1(n6628), .C2(keyinput36), 
        .A(n6627), .ZN(n6630) );
  NOR4_X1 U7534 ( .A1(n6633), .A2(n6632), .A3(n6631), .A4(n6630), .ZN(n6634)
         );
  NAND4_X1 U7535 ( .A1(n6637), .A2(n6636), .A3(n6635), .A4(n6634), .ZN(n6638)
         );
  NOR2_X1 U7536 ( .A1(n6639), .A2(n6638), .ZN(n6667) );
  NAND4_X1 U7537 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(
        INSTQUEUE_REG_13__3__SCAN_IN), .A3(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .A4(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6643) );
  NAND4_X1 U7538 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(
        INSTQUEUE_REG_9__6__SCAN_IN), .A3(PHYADDRPOINTER_REG_14__SCAN_IN), 
        .A4(DATAO_REG_23__SCAN_IN), .ZN(n6642) );
  NAND4_X1 U7539 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(
        INSTQUEUE_REG_14__3__SCAN_IN), .A3(REIP_REG_15__SCAN_IN), .A4(
        LWORD_REG_14__SCAN_IN), .ZN(n6641) );
  NAND4_X1 U7540 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A3(ADDRESS_REG_8__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6640) );
  NOR4_X1 U7541 ( .A1(n6643), .A2(n6642), .A3(n6641), .A4(n6640), .ZN(n6660)
         );
  NOR4_X1 U7542 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(
        STATE_REG_2__SCAN_IN), .A3(EBX_REG_9__SCAN_IN), .A4(EAX_REG_3__SCAN_IN), .ZN(n6647) );
  NOR4_X1 U7543 ( .A1(READY_N), .A2(EAX_REG_5__SCAN_IN), .A3(
        EAX_REG_6__SCAN_IN), .A4(LWORD_REG_6__SCAN_IN), .ZN(n6646) );
  NOR4_X1 U7544 ( .A1(STATE2_REG_0__SCAN_IN), .A2(DATAO_REG_29__SCAN_IN), .A3(
        DATAO_REG_24__SCAN_IN), .A4(LWORD_REG_7__SCAN_IN), .ZN(n6645) );
  NOR4_X1 U7545 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(EBX_REG_4__SCAN_IN), 
        .A3(EBX_REG_5__SCAN_IN), .A4(DATAI_0_), .ZN(n6644) );
  NAND4_X1 U7546 ( .A1(n6647), .A2(n6646), .A3(n6645), .A4(n6644), .ZN(n6653)
         );
  NAND4_X1 U7547 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        REIP_REG_3__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        ADDRESS_REG_19__SCAN_IN), .ZN(n6652) );
  NOR4_X1 U7548 ( .A1(EBX_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A3(REIP_REG_7__SCAN_IN), .A4(
        D_C_N_REG_SCAN_IN), .ZN(n6650) );
  NOR4_X1 U7549 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(
        INSTQUEUE_REG_13__4__SCAN_IN), .A3(INSTQUEUE_REG_7__2__SCAN_IN), .A4(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n6649) );
  NOR4_X1 U7550 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(
        INSTQUEUE_REG_8__4__SCAN_IN), .A3(EAX_REG_22__SCAN_IN), .A4(DATAI_30_), 
        .ZN(n6648) );
  NAND3_X1 U7551 ( .A1(n6650), .A2(n6649), .A3(n6648), .ZN(n6651) );
  NOR3_X1 U7552 ( .A1(n6653), .A2(n6652), .A3(n6651), .ZN(n6659) );
  NAND4_X1 U7553 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A3(DATAI_14_), .A4(DATAI_2_), .ZN(
        n6657) );
  NAND4_X1 U7554 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        EBX_REG_16__SCAN_IN), .A3(EAX_REG_17__SCAN_IN), .A4(
        PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6656) );
  NAND4_X1 U7555 ( .A1(EBX_REG_17__SCAN_IN), .A2(DATAI_3_), .A3(
        UWORD_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_26__SCAN_IN), .ZN(n6655) );
  NAND4_X1 U7556 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        EAX_REG_28__SCAN_IN), .A3(LWORD_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_4__SCAN_IN), .ZN(n6654) );
  NOR4_X1 U7557 ( .A1(n6657), .A2(n6656), .A3(n6655), .A4(n6654), .ZN(n6658)
         );
  NAND3_X1 U7558 ( .A1(n6660), .A2(n6659), .A3(n6658), .ZN(n6665) );
  AOI222_X1 U7559 ( .A1(n6663), .A2(ADDRESS_REG_5__SCAN_IN), .B1(
        REIP_REG_6__SCAN_IN), .B2(n6662), .C1(REIP_REG_7__SCAN_IN), .C2(n6661), 
        .ZN(n6664) );
  XNOR2_X1 U7560 ( .A(n6665), .B(n6664), .ZN(n6666) );
  XNOR2_X1 U7561 ( .A(n6667), .B(n6666), .ZN(U3189) );
  AND2_X2 U34470 ( .A1(n2959), .A2(n2960), .ZN(n3331) );
  AND4_X1 U4008 ( .A1(n3174), .A2(n3173), .A3(n3172), .A4(n3171), .ZN(n4262)
         );
  CLKBUF_X1 U3405 ( .A(n3935), .Z(n3822) );
  AOI22_X1 U3406 ( .A1(n6567), .A2(keyinput48), .B1(keyinput18), .B2(n6566), 
        .ZN(n6565) );
  CLKBUF_X1 U3454 ( .A(n4346), .Z(n4614) );
  NAND2_X1 U3467 ( .A1(n4153), .A2(n3458), .ZN(n4259) );
  CLKBUF_X1 U3553 ( .A(n3331), .Z(n3934) );
endmodule

