

module b14_C_gen_AntiSAT_k_256_1 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099;

  INV_X1 U2475 ( .A(n2564), .ZN(n2598) );
  CLKBUF_X2 U2476 ( .A(n2887), .Z(n2600) );
  INV_X2 U2477 ( .A(n2234), .ZN(n2917) );
  INV_X1 U2478 ( .A(n2945), .ZN(n2899) );
  INV_X1 U2479 ( .A(n2933), .ZN(n2913) );
  CLKBUF_X2 U2480 ( .A(n2948), .Z(n2234) );
  AND2_X1 U2483 ( .A1(n2479), .A2(n2478), .ZN(n2546) );
  NAND2_X1 U2484 ( .A1(n2311), .A2(IR_REG_31__SCAN_IN), .ZN(n3095) );
  OAI21_X1 U2485 ( .B1(n3111), .B2(n4710), .A(n2267), .ZN(n3108) );
  NAND2_X2 U2486 ( .A1(n2280), .A2(n2536), .ZN(n2770) );
  XNOR2_X2 U2487 ( .A(n2472), .B(IR_REG_30__SCAN_IN), .ZN(n3127) );
  NAND2_X1 U2488 ( .A1(n2507), .A2(n2981), .ZN(n2948) );
  AOI21_X1 U2489 ( .B1(n4283), .B2(n2357), .A(n2354), .ZN(n2353) );
  OR2_X1 U2490 ( .A1(n3669), .A2(n3670), .ZN(n3671) );
  NAND2_X1 U2491 ( .A1(n3747), .A2(n3746), .ZN(n3745) );
  NAND2_X1 U2492 ( .A1(n3936), .A2(n3939), .ZN(n3057) );
  INV_X2 U2493 ( .A(n4659), .ZN(n4658) );
  INV_X4 U2494 ( .A(n2770), .ZN(n2984) );
  INV_X1 U2495 ( .A(n2574), .ZN(n3017) );
  NAND4_X1 U2496 ( .A1(n2604), .A2(n2603), .A3(n2602), .A4(n2601), .ZN(n4069)
         );
  NAND3_X1 U2497 ( .A1(n2570), .A2(n2569), .A3(n2568), .ZN(n2574) );
  INV_X1 U2498 ( .A(n2553), .ZN(n2945) );
  INV_X1 U2499 ( .A(n3329), .ZN(n3331) );
  INV_X1 U2500 ( .A(n2507), .ZN(n2280) );
  AND2_X1 U2501 ( .A1(n2536), .A2(n2507), .ZN(n2553) );
  CLKBUF_X3 U2502 ( .A(n2565), .Z(n2840) );
  INV_X1 U2503 ( .A(n2996), .ZN(n4539) );
  NAND2_X1 U2504 ( .A1(n2528), .A2(IR_REG_31__SCAN_IN), .ZN(n2499) );
  NAND2_X1 U2505 ( .A1(n2503), .A2(n2502), .ZN(n2996) );
  INV_X1 U2506 ( .A(n3127), .ZN(n2478) );
  INV_X1 U2507 ( .A(n3241), .ZN(n3286) );
  BUF_X4 U2508 ( .A(n2552), .Z(n3133) );
  INV_X1 U2509 ( .A(n3118), .ZN(n2969) );
  NAND2_X1 U2510 ( .A1(n2471), .A2(IR_REG_31__SCAN_IN), .ZN(n2472) );
  AND2_X1 U2511 ( .A1(n2470), .A2(n2471), .ZN(n4538) );
  XNOR2_X1 U2512 ( .A(n2490), .B(IR_REG_26__SCAN_IN), .ZN(n3118) );
  MUX2_X1 U2513 ( .A(IR_REG_31__SCAN_IN), .B(n2469), .S(IR_REG_29__SCAN_IN), 
        .Z(n2470) );
  NOR2_X2 U2514 ( .A1(n2797), .A2(IR_REG_17__SCAN_IN), .ZN(n2800) );
  NAND2_X1 U2515 ( .A1(n2520), .A2(n2239), .ZN(n2797) );
  AND2_X1 U2516 ( .A1(n2308), .A2(n2374), .ZN(n2491) );
  AND2_X1 U2517 ( .A1(n4999), .A2(n2461), .ZN(n2426) );
  INV_X1 U2518 ( .A(IR_REG_25__SCAN_IN), .ZN(n2466) );
  INV_X1 U2519 ( .A(IR_REG_20__SCAN_IN), .ZN(n2498) );
  NOR2_X1 U2520 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2459)
         );
  NOR2_X1 U2521 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2457)
         );
  INV_X1 U2522 ( .A(IR_REG_3__SCAN_IN), .ZN(n2586) );
  INV_X1 U2523 ( .A(IR_REG_13__SCAN_IN), .ZN(n2461) );
  NOR2_X1 U2524 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2458)
         );
  INV_X2 U2525 ( .A(IR_REG_14__SCAN_IN), .ZN(n4999) );
  NOR2_X1 U2526 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2462)
         );
  NOR2_X1 U2527 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2484)
         );
  NAND2_X1 U2528 ( .A1(n3311), .A2(n2506), .ZN(n4694) );
  OAI21_X2 U2529 ( .B1(n3522), .B2(n3034), .A(n3033), .ZN(n3571) );
  OAI22_X2 U2530 ( .A1(n3489), .A2(n3032), .B1(n3502), .B2(n3546), .ZN(n3522)
         );
  OR2_X1 U2531 ( .A1(n4192), .A2(n4211), .ZN(n3051) );
  INV_X1 U2532 ( .A(n2272), .ZN(n2271) );
  OAI21_X1 U2533 ( .B1(n2497), .B2(n2761), .A(n4826), .ZN(n2272) );
  NAND2_X1 U2534 ( .A1(n2428), .A2(n2429), .ZN(n2787) );
  AOI21_X1 U2535 ( .B1(n2431), .B2(n2435), .A(n2430), .ZN(n2429) );
  INV_X1 U2536 ( .A(n3651), .ZN(n2430) );
  NOR2_X1 U2537 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2464)
         );
  NOR2_X1 U2538 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2463)
         );
  AND2_X1 U2539 ( .A1(n2239), .A2(n2243), .ZN(n2308) );
  AND2_X1 U2540 ( .A1(n2467), .A2(n2466), .ZN(n2437) );
  INV_X1 U2541 ( .A(IR_REG_26__SCAN_IN), .ZN(n2467) );
  OR2_X1 U2542 ( .A1(n2753), .A2(n2435), .ZN(n2433) );
  NAND2_X1 U2543 ( .A1(n3259), .A2(n3258), .ZN(n2414) );
  XNOR2_X1 U2544 ( .A(n2573), .B(n2917), .ZN(n2578) );
  XNOR2_X1 U2545 ( .A(n3453), .B(n4665), .ZN(n4588) );
  INV_X1 U2546 ( .A(n2375), .ZN(n2283) );
  OAI22_X1 U2547 ( .A1(n4118), .A2(n4117), .B1(REG2_REG_13__SCAN_IN), .B2(
        n4541), .ZN(n4119) );
  NOR2_X1 U2548 ( .A1(n4029), .A2(n3090), .ZN(n4161) );
  NOR2_X1 U2549 ( .A1(n2885), .A2(n4975), .ZN(n2907) );
  NOR2_X1 U2550 ( .A1(n4212), .A2(n4237), .ZN(n3049) );
  AOI21_X1 U2551 ( .B1(n2339), .B2(n3920), .A(n2249), .ZN(n2341) );
  AND2_X1 U2552 ( .A1(n4038), .A2(n3092), .ZN(n4334) );
  NAND2_X1 U2553 ( .A1(n2496), .A2(n2953), .ZN(n2536) );
  INV_X1 U2554 ( .A(n4540), .ZN(n4144) );
  XNOR2_X1 U2555 ( .A(n2379), .B(n4141), .ZN(n2378) );
  NAND2_X1 U2556 ( .A1(n2381), .A2(n2380), .ZN(n2379) );
  NAND2_X1 U2557 ( .A1(n4138), .A2(REG1_REG_18__SCAN_IN), .ZN(n2380) );
  NOR2_X1 U2558 ( .A1(n3808), .A2(n3807), .ZN(n2435) );
  NAND2_X1 U2559 ( .A1(n2410), .A2(n3745), .ZN(n2275) );
  AND2_X1 U2560 ( .A1(n2406), .A2(n3635), .ZN(n2405) );
  INV_X1 U2561 ( .A(n2945), .ZN(n2914) );
  INV_X1 U2562 ( .A(n4538), .ZN(n2479) );
  OAI21_X1 U2563 ( .B1(n3220), .B2(n2263), .A(n2382), .ZN(n3164) );
  NAND2_X1 U2564 ( .A1(n4543), .A2(REG1_REG_7__SCAN_IN), .ZN(n2382) );
  AND2_X1 U2565 ( .A1(n4185), .A2(n4407), .ZN(n4028) );
  INV_X1 U2566 ( .A(n2295), .ZN(n2294) );
  AND2_X1 U2567 ( .A1(n2298), .A2(n4022), .ZN(n2295) );
  NOR2_X1 U2568 ( .A1(n2301), .A2(n2300), .ZN(n2299) );
  INV_X1 U2569 ( .A(n2304), .ZN(n2300) );
  OR2_X1 U2570 ( .A1(n2302), .A2(n2301), .ZN(n2298) );
  NOR2_X1 U2571 ( .A1(n2306), .A2(n2305), .ZN(n2304) );
  INV_X1 U2572 ( .A(n4019), .ZN(n2305) );
  INV_X1 U2573 ( .A(n2256), .ZN(n2306) );
  NAND2_X1 U2574 ( .A1(n2303), .A2(n2256), .ZN(n2302) );
  INV_X1 U2575 ( .A(n4024), .ZN(n2303) );
  NOR2_X1 U2576 ( .A1(n2352), .A2(n2349), .ZN(n2348) );
  INV_X1 U2577 ( .A(n3043), .ZN(n2352) );
  INV_X1 U2578 ( .A(n4348), .ZN(n2349) );
  NAND2_X1 U2579 ( .A1(n2351), .A2(n3043), .ZN(n2350) );
  INV_X1 U2580 ( .A(n3041), .ZN(n2351) );
  OR2_X1 U2581 ( .A1(n4366), .A2(n4245), .ZN(n4325) );
  AOI21_X1 U2582 ( .B1(n3075), .B2(n3906), .A(n2289), .ZN(n2288) );
  INV_X1 U2583 ( .A(n3958), .ZN(n2289) );
  INV_X1 U2584 ( .A(n3075), .ZN(n2290) );
  NOR2_X1 U2585 ( .A1(n3872), .A2(n4211), .ZN(n2322) );
  NOR2_X1 U2586 ( .A1(n4296), .A2(n4306), .ZN(n2316) );
  INV_X1 U2587 ( .A(n3656), .ZN(n3581) );
  INV_X1 U2588 ( .A(IR_REG_15__SCAN_IN), .ZN(n4996) );
  INV_X1 U2589 ( .A(IR_REG_2__SCAN_IN), .ZN(n2279) );
  AND2_X1 U2590 ( .A1(n2407), .A2(n2409), .ZN(n2410) );
  NAND2_X1 U2591 ( .A1(n3808), .A2(n3807), .ZN(n2434) );
  OR2_X1 U2592 ( .A1(n2873), .A2(n2872), .ZN(n2885) );
  AOI21_X1 U2593 ( .B1(n2424), .B2(n2422), .A(n2265), .ZN(n2421) );
  NAND2_X1 U2594 ( .A1(n2401), .A2(n3765), .ZN(n3730) );
  OR2_X1 U2595 ( .A1(n3767), .A2(n3768), .ZN(n2401) );
  OAI21_X1 U2596 ( .B1(n3820), .B2(n2396), .A(n2395), .ZN(n3765) );
  NAND2_X1 U2597 ( .A1(n2240), .A2(n2397), .ZN(n2396) );
  AOI21_X1 U2598 ( .B1(n2402), .B2(n2240), .A(n2261), .ZN(n2395) );
  INV_X1 U2599 ( .A(n3821), .ZN(n2397) );
  OAI21_X1 U2600 ( .B1(n3820), .B2(n2400), .A(n2398), .ZN(n3767) );
  OR2_X1 U2601 ( .A1(n2892), .A2(n3821), .ZN(n2400) );
  OR2_X1 U2602 ( .A1(n2399), .A2(n2892), .ZN(n2398) );
  NAND2_X1 U2603 ( .A1(n2240), .A2(n2261), .ZN(n2892) );
  NAND2_X1 U2604 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2512) );
  NOR2_X1 U2605 ( .A1(n2731), .A2(n2730), .ZN(n2733) );
  NAND2_X1 U2606 ( .A1(n2752), .A2(n2751), .ZN(n2753) );
  NAND2_X1 U2607 ( .A1(n3671), .A2(n2250), .ZN(n2752) );
  INV_X1 U2608 ( .A(n3797), .ZN(n2861) );
  NAND2_X1 U2609 ( .A1(n2849), .A2(REG3_REG_21__SCAN_IN), .ZN(n2873) );
  INV_X1 U2610 ( .A(n3251), .ZN(n2281) );
  OR2_X1 U2611 ( .A1(n2564), .A2(n2530), .ZN(n2531) );
  XNOR2_X1 U2612 ( .A(n3142), .B(n4547), .ZN(n4096) );
  NOR2_X1 U2613 ( .A1(n3179), .A2(n2329), .ZN(n2328) );
  NOR2_X1 U2614 ( .A1(n3179), .A2(n3214), .ZN(n2327) );
  INV_X1 U2615 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2329) );
  AND2_X1 U2616 ( .A1(n2331), .A2(n2330), .ZN(n3166) );
  NAND2_X1 U2617 ( .A1(n4545), .A2(REG2_REG_5__SCAN_IN), .ZN(n2330) );
  NOR2_X1 U2618 ( .A1(n3163), .A2(n2383), .ZN(n3220) );
  NOR2_X1 U2619 ( .A1(n3162), .A2(n2384), .ZN(n2383) );
  INV_X1 U2620 ( .A(n4544), .ZN(n2384) );
  AOI21_X1 U2621 ( .B1(n4123), .B2(REG2_REG_15__SCAN_IN), .A(n2248), .ZN(n4125) );
  NAND2_X1 U2622 ( .A1(n4609), .A2(n4107), .ZN(n4108) );
  NAND2_X1 U2623 ( .A1(n2262), .A2(n2241), .ZN(n2370) );
  INV_X1 U2624 ( .A(n4193), .ZN(n2373) );
  OAI21_X1 U2625 ( .B1(n2356), .B2(n3045), .A(n2447), .ZN(n2354) );
  NOR2_X1 U2626 ( .A1(n4283), .A2(n2361), .ZN(n2359) );
  OR2_X1 U2627 ( .A1(n4370), .A2(n4349), .ZN(n3041) );
  AND2_X1 U2628 ( .A1(n4056), .A2(n4383), .ZN(n3038) );
  NAND2_X1 U2629 ( .A1(n4345), .A2(n4348), .ZN(n4344) );
  NOR2_X1 U2630 ( .A1(n2255), .A2(n2377), .ZN(n2376) );
  NAND2_X1 U2631 ( .A1(n3571), .A2(n3906), .ZN(n3570) );
  NOR2_X1 U2632 ( .A1(n3025), .A2(n2338), .ZN(n2345) );
  INV_X1 U2633 ( .A(n3023), .ZN(n2338) );
  OAI21_X1 U2634 ( .B1(n3025), .B2(n2340), .A(n2254), .ZN(n2339) );
  NAND2_X1 U2635 ( .A1(n3023), .A2(n3024), .ZN(n2340) );
  OAI21_X1 U2636 ( .B1(n3300), .B2(n3060), .A(n3945), .ZN(n3340) );
  INV_X1 U2637 ( .A(n4369), .ZN(n4331) );
  NAND2_X1 U2638 ( .A1(n3286), .A2(n3310), .ZN(n3329) );
  AND2_X1 U2639 ( .A1(n4197), .A2(n4170), .ZN(n4172) );
  NOR2_X1 U2640 ( .A1(n4233), .A2(n2319), .ZN(n4197) );
  INV_X1 U2641 ( .A(n2322), .ZN(n2319) );
  OR2_X1 U2642 ( .A1(n4262), .A2(n4237), .ZN(n4233) );
  INV_X1 U2643 ( .A(n4054), .ZN(n4425) );
  INV_X1 U2644 ( .A(n4059), .ZN(n3595) );
  AND2_X1 U2645 ( .A1(n4312), .A2(n4674), .ZN(n4468) );
  AND2_X1 U2646 ( .A1(n3148), .A2(n3131), .ZN(n4408) );
  NAND2_X1 U2647 ( .A1(n2955), .A2(n3118), .ZN(n3136) );
  INV_X1 U2648 ( .A(IR_REG_29__SCAN_IN), .ZN(n4797) );
  NAND3_X1 U2649 ( .A1(n2246), .A2(n2308), .A3(n2374), .ZN(n2468) );
  NAND2_X1 U2650 ( .A1(n2394), .A2(IR_REG_31__SCAN_IN), .ZN(n2393) );
  INV_X1 U2651 ( .A(IR_REG_23__SCAN_IN), .ZN(n2970) );
  AND2_X1 U2652 ( .A1(n2970), .A2(IR_REG_24__SCAN_IN), .ZN(n2392) );
  NAND2_X1 U2653 ( .A1(n2488), .A2(IR_REG_31__SCAN_IN), .ZN(n2971) );
  NOR2_X1 U2654 ( .A1(n2441), .A2(IR_REG_22__SCAN_IN), .ZN(n2440) );
  XNOR2_X1 U2655 ( .A(n2971), .B(n2970), .ZN(n3132) );
  NOR2_X1 U2656 ( .A1(n2689), .A2(IR_REG_9__SCAN_IN), .ZN(n2721) );
  INV_X1 U2657 ( .A(IR_REG_7__SCAN_IN), .ZN(n4798) );
  AND2_X1 U2658 ( .A1(n2937), .A2(n2926), .ZN(n4173) );
  AND2_X1 U2659 ( .A1(n3007), .A2(n2974), .ZN(n3883) );
  INV_X1 U2660 ( .A(n4273), .ZN(n4308) );
  OAI21_X1 U2661 ( .B1(n4200), .B2(n2284), .A(n2912), .ZN(n4409) );
  NAND2_X1 U2662 ( .A1(n2898), .A2(n2897), .ZN(n4192) );
  XNOR2_X1 U2663 ( .A(n3166), .B(n4544), .ZN(n3168) );
  NAND2_X1 U2664 ( .A1(n4586), .A2(n3454), .ZN(n4118) );
  XNOR2_X1 U2665 ( .A(n4119), .B(n2336), .ZN(n4597) );
  NOR2_X1 U2666 ( .A1(n4597), .A2(n4598), .ZN(n4596) );
  XNOR2_X1 U2667 ( .A(n4108), .B(n4124), .ZN(n4618) );
  NOR2_X1 U2668 ( .A1(n4618), .A2(REG1_REG_16__SCAN_IN), .ZN(n4619) );
  NOR2_X1 U2669 ( .A1(n4128), .A2(n4129), .ZN(n4135) );
  AND2_X1 U2670 ( .A1(n4077), .A2(n4074), .ZN(n4629) );
  OR2_X1 U2671 ( .A1(n4135), .A2(n2333), .ZN(n2332) );
  AND2_X1 U2672 ( .A1(n4138), .A2(REG2_REG_18__SCAN_IN), .ZN(n2333) );
  INV_X1 U2673 ( .A(n4587), .ZN(n4622) );
  INV_X1 U2674 ( .A(n2366), .ZN(n2365) );
  AND2_X1 U2675 ( .A1(n2528), .A2(n2527), .ZN(n4540) );
  NAND2_X1 U2676 ( .A1(n2270), .A2(IR_REG_31__SCAN_IN), .ZN(n2526) );
  NOR2_X1 U2677 ( .A1(n2432), .A2(n3650), .ZN(n2431) );
  INV_X1 U2678 ( .A(n2434), .ZN(n2432) );
  NOR2_X1 U2679 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2460)
         );
  AND2_X1 U2680 ( .A1(n2486), .A2(n2444), .ZN(n2443) );
  INV_X1 U2681 ( .A(IR_REG_17__SCAN_IN), .ZN(n2444) );
  INV_X1 U2682 ( .A(IR_REG_10__SCAN_IN), .ZN(n5001) );
  NAND2_X1 U2683 ( .A1(n2412), .A2(n3856), .ZN(n2409) );
  NAND2_X1 U2684 ( .A1(n2633), .A2(n2413), .ZN(n2412) );
  NAND2_X1 U2685 ( .A1(n3855), .A2(n2408), .ZN(n2407) );
  INV_X1 U2686 ( .A(n2633), .ZN(n2408) );
  INV_X1 U2687 ( .A(n2402), .ZN(n2399) );
  INV_X1 U2688 ( .A(IR_REG_27__SCAN_IN), .ZN(n4799) );
  INV_X1 U2689 ( .A(n2714), .ZN(n2427) );
  INV_X1 U2690 ( .A(n2920), .ZN(n2947) );
  CLKBUF_X1 U2691 ( .A(n2933), .Z(n2946) );
  AND2_X1 U2692 ( .A1(n3912), .A2(n4227), .ZN(n4024) );
  NAND2_X1 U2693 ( .A1(n4548), .A2(REG2_REG_2__SCAN_IN), .ZN(n2326) );
  NOR2_X1 U2694 ( .A1(n3198), .A2(n2325), .ZN(n3142) );
  INV_X1 U2695 ( .A(n2326), .ZN(n2325) );
  AND2_X1 U2696 ( .A1(n4302), .A2(n3080), .ZN(n4249) );
  OR2_X1 U2697 ( .A1(n4325), .A2(n4247), .ZN(n4303) );
  INV_X1 U2698 ( .A(n3035), .ZN(n2377) );
  NAND2_X1 U2699 ( .A1(n4011), .A2(n3573), .ZN(n3572) );
  AND2_X1 U2700 ( .A1(n2345), .A2(n3920), .ZN(n2337) );
  NAND2_X1 U2701 ( .A1(n3385), .A2(n3781), .ZN(n3942) );
  NAND2_X1 U2702 ( .A1(n4070), .A2(n3286), .ZN(n3932) );
  AND2_X1 U2703 ( .A1(n3508), .A2(n3546), .ZN(n2313) );
  OR2_X1 U2704 ( .A1(n3136), .A2(D_REG_1__SCAN_IN), .ZN(n3100) );
  NAND2_X1 U2705 ( .A1(n2443), .A2(n2442), .ZN(n2441) );
  INV_X1 U2706 ( .A(IR_REG_21__SCAN_IN), .ZN(n2442) );
  OR2_X1 U2707 ( .A1(n2797), .A2(n2439), .ZN(n2500) );
  INV_X1 U2708 ( .A(n2443), .ZN(n2439) );
  NOR2_X1 U2709 ( .A1(n2797), .A2(n2441), .ZN(n2504) );
  XNOR2_X1 U2710 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_f56), .ZN(n5034) );
  INV_X1 U2711 ( .A(IR_REG_6__SCAN_IN), .ZN(n5011) );
  XNOR2_X1 U2712 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_g56), .ZN(n4829) );
  NOR2_X1 U2713 ( .A1(n3856), .A2(n3855), .ZN(n2411) );
  NAND2_X1 U2714 ( .A1(n2404), .A2(n2403), .ZN(n2402) );
  INV_X1 U2715 ( .A(n3663), .ZN(n2403) );
  INV_X1 U2716 ( .A(n3662), .ZN(n2404) );
  XNOR2_X1 U2717 ( .A(n2591), .B(n2234), .ZN(n2594) );
  NAND2_X1 U2718 ( .A1(n2421), .A2(n2419), .ZN(n2418) );
  NAND2_X1 U2719 ( .A1(n2952), .A2(n2423), .ZN(n2419) );
  NAND2_X1 U2720 ( .A1(n2405), .A2(n2275), .ZN(n2274) );
  NAND2_X1 U2721 ( .A1(n3879), .A2(n3881), .ZN(n2276) );
  NOR2_X1 U2722 ( .A1(n3878), .A2(n3737), .ZN(n2277) );
  CLKBUF_X1 U2723 ( .A(n3701), .Z(n3800) );
  AND2_X1 U2724 ( .A1(n2552), .A2(DATAI_22_), .ZN(n3046) );
  NAND2_X1 U2725 ( .A1(n3671), .A2(n2714), .ZN(n3834) );
  INV_X1 U2726 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3850) );
  AND2_X1 U2727 ( .A1(n2617), .A2(REG3_REG_5__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U2728 ( .A1(n2755), .A2(n2476), .ZN(n2772) );
  AND3_X1 U2729 ( .A1(n3109), .A2(n3279), .A3(n3100), .ZN(n3007) );
  OAI21_X1 U2730 ( .B1(n4548), .B2(REG2_REG_2__SCAN_IN), .A(n2326), .ZN(n3200)
         );
  AOI21_X1 U2731 ( .B1(n4083), .B2(n3199), .A(n3200), .ZN(n3198) );
  NAND2_X1 U2732 ( .A1(n3211), .A2(REG1_REG_4__SCAN_IN), .ZN(n3210) );
  INV_X1 U2733 ( .A(n3164), .ZN(n3429) );
  NAND2_X1 U2734 ( .A1(n4578), .A2(n3451), .ZN(n3453) );
  NAND2_X1 U2735 ( .A1(n4588), .A2(REG2_REG_12__SCAN_IN), .ZN(n4586) );
  AND2_X1 U2736 ( .A1(n3134), .A2(n3133), .ZN(n3146) );
  NOR2_X1 U2737 ( .A1(n4632), .A2(n4110), .ZN(n4140) );
  NAND2_X1 U2738 ( .A1(n4140), .A2(n4139), .ZN(n2381) );
  NOR2_X1 U2739 ( .A1(n4161), .A2(n2369), .ZN(n2368) );
  INV_X1 U2740 ( .A(n2370), .ZN(n2369) );
  OAI22_X1 U2741 ( .A1(n4161), .A2(n2367), .B1(n4157), .B2(n3624), .ZN(n2366)
         );
  NAND2_X1 U2742 ( .A1(n2370), .A2(n2372), .ZN(n2367) );
  OR2_X1 U2743 ( .A1(n4028), .A2(n3995), .ZN(n4177) );
  AOI21_X1 U2744 ( .B1(n2295), .B2(n2293), .A(n3993), .ZN(n2292) );
  INV_X1 U2745 ( .A(n2299), .ZN(n2293) );
  NAND2_X1 U2746 ( .A1(n2296), .A2(n2298), .ZN(n4187) );
  NAND2_X1 U2747 ( .A1(n3088), .A2(n2299), .ZN(n2296) );
  OR2_X1 U2748 ( .A1(n3900), .A2(n3993), .ZN(n4195) );
  NAND2_X1 U2749 ( .A1(n2297), .A2(n2302), .ZN(n4209) );
  NAND2_X1 U2750 ( .A1(n3088), .A2(n2304), .ZN(n2297) );
  AOI21_X1 U2751 ( .B1(n4243), .B2(n3048), .A(n3047), .ZN(n4226) );
  AND2_X1 U2752 ( .A1(n4054), .A2(n4260), .ZN(n3047) );
  NAND2_X1 U2753 ( .A1(n2552), .A2(DATAI_23_), .ZN(n4254) );
  AND2_X1 U2754 ( .A1(n4284), .A2(n4250), .ZN(n4270) );
  AND4_X1 U2755 ( .A1(n2866), .A2(n2865), .A3(n2864), .A4(n2863), .ZN(n4288)
         );
  AND2_X1 U2756 ( .A1(n3901), .A2(n4250), .ZN(n4285) );
  NAND2_X1 U2757 ( .A1(n2347), .A2(n2260), .ZN(n4301) );
  AND2_X1 U2758 ( .A1(n2838), .A2(n2837), .ZN(n2849) );
  NOR2_X1 U2759 ( .A1(n2808), .A2(n3850), .ZN(n2838) );
  INV_X1 U2760 ( .A(n4349), .ZN(n4357) );
  AOI21_X1 U2761 ( .B1(n2288), .B2(n2290), .A(n3613), .ZN(n2287) );
  NAND2_X1 U2762 ( .A1(n2286), .A2(n2288), .ZN(n3614) );
  OR2_X1 U2763 ( .A1(n4011), .A2(n2290), .ZN(n2286) );
  AND2_X1 U2764 ( .A1(n2733), .A2(REG3_REG_13__SCAN_IN), .ZN(n2755) );
  OAI21_X1 U2765 ( .B1(n3532), .B2(n3029), .A(n3028), .ZN(n3501) );
  OAI21_X1 U2766 ( .B1(n3412), .B2(n3969), .A(n3952), .ZN(n3533) );
  NOR2_X1 U2767 ( .A1(n2679), .A2(n2473), .ZN(n2699) );
  NAND2_X1 U2768 ( .A1(n2307), .A2(n3950), .ZN(n3412) );
  NAND2_X1 U2769 ( .A1(n3473), .A2(n3953), .ZN(n2307) );
  INV_X1 U2770 ( .A(n3638), .ZN(n3360) );
  OAI21_X1 U2771 ( .B1(n3340), .B2(n3338), .A(n3961), .ZN(n3367) );
  NAND2_X1 U2772 ( .A1(n3059), .A2(n3941), .ZN(n3300) );
  INV_X1 U2773 ( .A(n4334), .ZN(n4367) );
  OAI21_X1 U2774 ( .B1(n3056), .B2(n3931), .A(n3935), .ZN(n3318) );
  INV_X1 U2775 ( .A(n3312), .ZN(n3310) );
  AND2_X1 U2776 ( .A1(n3189), .A2(n3131), .ZN(n4369) );
  INV_X1 U2777 ( .A(n2975), .ZN(n3311) );
  AND2_X1 U2778 ( .A1(n3103), .A2(n3137), .ZN(n3279) );
  NAND2_X1 U2779 ( .A1(n2536), .A2(n4660), .ZN(n3275) );
  NOR2_X1 U2780 ( .A1(n4394), .A2(n4395), .ZN(n4393) );
  INV_X1 U2781 ( .A(n4148), .ZN(n4395) );
  NAND2_X1 U2782 ( .A1(n2323), .A2(n2322), .ZN(n2321) );
  NOR2_X1 U2783 ( .A1(n4407), .A2(n2324), .ZN(n2323) );
  OR2_X1 U2784 ( .A1(n4156), .A2(n4000), .ZN(n4394) );
  NAND2_X1 U2785 ( .A1(n2552), .A2(DATAI_25_), .ZN(n4219) );
  NOR2_X1 U2786 ( .A1(n4233), .A2(n4211), .ZN(n4217) );
  NAND2_X1 U2787 ( .A1(n2316), .A2(n4276), .ZN(n2315) );
  NOR2_X1 U2788 ( .A1(n4338), .A2(n2314), .ZN(n4291) );
  INV_X1 U2789 ( .A(n2316), .ZN(n2314) );
  INV_X1 U2790 ( .A(n4296), .ZN(n4440) );
  AND2_X1 U2791 ( .A1(n4374), .A2(n4357), .ZN(n4355) );
  NAND2_X1 U2792 ( .A1(n4355), .A2(n4336), .ZN(n4338) );
  NOR2_X1 U2793 ( .A1(n4373), .A2(n4383), .ZN(n4374) );
  OR2_X1 U2794 ( .A1(n3607), .A2(n3739), .ZN(n4373) );
  OR2_X1 U2795 ( .A1(n4476), .A2(n3888), .ZN(n3607) );
  NAND2_X1 U2796 ( .A1(n2238), .A2(n3581), .ZN(n4476) );
  NAND2_X1 U2797 ( .A1(n3529), .A2(n2313), .ZN(n3523) );
  NAND2_X1 U2798 ( .A1(n3529), .A2(n3508), .ZN(n3507) );
  INV_X1 U2799 ( .A(n3674), .ZN(n3534) );
  AND2_X1 U2800 ( .A1(n3531), .A2(n3534), .ZN(n3529) );
  NOR2_X1 U2801 ( .A1(n3470), .A2(n3790), .ZN(n3531) );
  OR2_X1 U2802 ( .A1(n3469), .A2(n3696), .ZN(n3470) );
  NOR2_X1 U2803 ( .A1(n3861), .A2(n3749), .ZN(n2312) );
  INV_X1 U2804 ( .A(n4459), .ZN(n4406) );
  NAND2_X1 U2805 ( .A1(n4678), .A2(n2237), .ZN(n3344) );
  NAND2_X1 U2806 ( .A1(n4678), .A2(n3395), .ZN(n3296) );
  INV_X1 U2807 ( .A(n4408), .ZN(n4460) );
  NAND2_X1 U2808 ( .A1(n2491), .A2(n2437), .ZN(n2311) );
  XNOR2_X1 U2809 ( .A(n2505), .B(n2487), .ZN(n2995) );
  OR2_X1 U2810 ( .A1(n2504), .A2(n2761), .ZN(n2505) );
  INV_X1 U2811 ( .A(IR_REG_19__SCAN_IN), .ZN(n4826) );
  INV_X1 U2812 ( .A(IR_REG_18__SCAN_IN), .ZN(n2497) );
  AND2_X1 U2813 ( .A1(n2778), .A2(n2510), .ZN(n4123) );
  INV_X1 U2814 ( .A(n2585), .ZN(n2456) );
  NAND2_X1 U2815 ( .A1(n2433), .A2(n2434), .ZN(n3654) );
  NAND2_X1 U2816 ( .A1(n3249), .A2(n2579), .ZN(n3259) );
  NAND2_X1 U2817 ( .A1(n2417), .A2(n2420), .ZN(n2416) );
  NAND2_X1 U2818 ( .A1(n2424), .A2(n2425), .ZN(n2420) );
  INV_X1 U2819 ( .A(n4219), .ZN(n4211) );
  INV_X1 U2820 ( .A(n4458), .ZN(n4383) );
  AND2_X1 U2821 ( .A1(n2552), .A2(DATAI_20_), .ZN(n4306) );
  INV_X1 U2822 ( .A(n3046), .ZN(n4276) );
  OR2_X1 U2823 ( .A1(n3702), .A2(n3703), .ZN(n2862) );
  NOR2_X1 U2824 ( .A1(n3701), .A2(n3796), .ZN(n2278) );
  NOR2_X1 U2825 ( .A1(n3820), .A2(n3821), .ZN(n3819) );
  NAND2_X1 U2826 ( .A1(n3745), .A2(n2633), .ZN(n3858) );
  NAND2_X2 U2827 ( .A1(n2987), .A2(n3232), .ZN(n3890) );
  NAND2_X1 U2828 ( .A1(n2840), .A2(REG2_REG_0__SCAN_IN), .ZN(n2535) );
  INV_X2 U2829 ( .A(U4043), .ZN(n4071) );
  NAND2_X1 U2830 ( .A1(n4084), .A2(n2236), .ZN(n4083) );
  AND2_X1 U2831 ( .A1(n3210), .A2(n2385), .ZN(n3177) );
  NAND2_X1 U2832 ( .A1(n3156), .A2(n4546), .ZN(n2385) );
  AOI21_X1 U2833 ( .B1(n3209), .B2(REG2_REG_4__SCAN_IN), .A(n2269), .ZN(n3180)
         );
  AOI22_X1 U2834 ( .A1(n3168), .A2(REG2_REG_6__SCAN_IN), .B1(n4544), .B2(n3167), .ZN(n3226) );
  AND2_X1 U2835 ( .A1(n4077), .A2(n3149), .ZN(n4587) );
  NOR2_X1 U2836 ( .A1(n4596), .A2(n4121), .ZN(n4606) );
  NOR2_X1 U2837 ( .A1(n4619), .A2(n4109), .ZN(n4631) );
  NAND2_X1 U2838 ( .A1(n4624), .A2(n2334), .ZN(n4128) );
  NAND2_X1 U2839 ( .A1(n4662), .A2(n2335), .ZN(n2334) );
  INV_X1 U2840 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2335) );
  NAND2_X1 U2841 ( .A1(n2364), .A2(n2370), .ZN(n4155) );
  NAND2_X1 U2842 ( .A1(n2373), .A2(n2371), .ZN(n2364) );
  AND2_X1 U2843 ( .A1(n2932), .A2(n2931), .ZN(n4185) );
  OR2_X1 U2844 ( .A1(n2925), .A2(n2908), .ZN(n4200) );
  NAND2_X1 U2845 ( .A1(n3088), .A2(n4019), .ZN(n4228) );
  INV_X1 U2846 ( .A(n2359), .ZN(n2355) );
  NAND2_X1 U2847 ( .A1(n4344), .A2(n3041), .ZN(n4323) );
  NAND2_X1 U2848 ( .A1(n3570), .A2(n3035), .ZN(n3557) );
  INV_X1 U2849 ( .A(n2339), .ZN(n2343) );
  NAND2_X1 U2850 ( .A1(n3337), .A2(n2345), .ZN(n2344) );
  OR2_X1 U2851 ( .A1(n3337), .A2(n3024), .ZN(n2346) );
  INV_X1 U2852 ( .A(n3262), .ZN(n3395) );
  NOR2_X1 U2853 ( .A1(n3329), .A2(n3106), .ZN(n4678) );
  NAND2_X1 U2854 ( .A1(n3233), .A2(n2997), .ZN(n4645) );
  INV_X1 U2855 ( .A(n3101), .ZN(n2997) );
  OR2_X1 U2856 ( .A1(n4360), .A2(n4694), .ZN(n4385) );
  OAI21_X1 U2857 ( .B1(n3622), .B2(n4468), .A(n2310), .ZN(n2309) );
  AOI21_X1 U2858 ( .B1(n4179), .B2(n4408), .A(n3099), .ZN(n2310) );
  OAI21_X1 U2859 ( .B1(n2320), .B2(n3107), .A(n4394), .ZN(n3627) );
  OR2_X1 U2860 ( .A1(n4172), .A2(n4171), .ZN(n4494) );
  OR2_X1 U2861 ( .A1(n3110), .A2(n3109), .ZN(n4700) );
  NAND2_X1 U2862 ( .A1(n3136), .A2(n3233), .ZN(n4659) );
  INV_X1 U2863 ( .A(n2468), .ZN(n2991) );
  INV_X1 U2864 ( .A(n2493), .ZN(n2495) );
  INV_X1 U2865 ( .A(n2390), .ZN(n2389) );
  NAND2_X1 U2866 ( .A1(n2971), .A2(n2392), .ZN(n2391) );
  OAI22_X1 U2867 ( .A1(n2393), .A2(n2970), .B1(IR_REG_31__SCAN_IN), .B2(n2394), 
        .ZN(n2390) );
  AND2_X1 U2868 ( .A1(n3132), .A2(STATE_REG_SCAN_IN), .ZN(n4660) );
  INV_X1 U2869 ( .A(n2995), .ZN(n4048) );
  XNOR2_X1 U2870 ( .A(n2815), .B(IR_REG_18__SCAN_IN), .ZN(n4138) );
  NOR2_X1 U2871 ( .A1(n2690), .A2(n2721), .ZN(n4553) );
  AND2_X1 U2872 ( .A1(n2668), .A2(n2655), .ZN(n4543) );
  AND2_X1 U2873 ( .A1(n2605), .A2(n2588), .ZN(n4547) );
  XNOR2_X1 U2874 ( .A(n2332), .B(n4136), .ZN(n4147) );
  AOI21_X1 U2875 ( .B1(n2378), .B2(n4629), .A(n4145), .ZN(n4146) );
  AND2_X1 U2876 ( .A1(n2586), .A2(n2455), .ZN(n2235) );
  AND2_X1 U2877 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2236)
         );
  AND2_X1 U2878 ( .A1(n3297), .A2(n3395), .ZN(n2237) );
  AND2_X1 U2879 ( .A1(n3529), .A2(n2259), .ZN(n2238) );
  AND2_X2 U2880 ( .A1(n2426), .A2(n2252), .ZN(n2239) );
  INV_X1 U2881 ( .A(n3861), .ZN(n3370) );
  NAND2_X1 U2882 ( .A1(n2355), .A2(n2357), .ZN(n4268) );
  NAND2_X1 U2883 ( .A1(n2520), .A2(n2426), .ZN(n2508) );
  OR2_X1 U2884 ( .A1(n2884), .A2(n2883), .ZN(n2240) );
  OR2_X1 U2885 ( .A1(n4185), .A2(n4170), .ZN(n2241) );
  INV_X1 U2886 ( .A(n3867), .ZN(n2422) );
  AND2_X1 U2887 ( .A1(n2417), .A2(n2266), .ZN(n2242) );
  INV_X2 U2888 ( .A(n4710), .ZN(n4713) );
  AND2_X1 U2889 ( .A1(n2552), .A2(DATAI_27_), .ZN(n4407) );
  INV_X1 U2890 ( .A(IR_REG_31__SCAN_IN), .ZN(n2761) );
  AND4_X1 U2891 ( .A1(n2458), .A2(n2459), .A3(n2460), .A4(n2457), .ZN(n2243)
         );
  OR2_X1 U2892 ( .A1(n4338), .A2(n2315), .ZN(n2244) );
  AND2_X1 U2893 ( .A1(n4799), .A2(n2437), .ZN(n2245) );
  AOI21_X1 U2894 ( .B1(n4226), .B2(n3050), .A(n3049), .ZN(n4206) );
  AND2_X1 U2895 ( .A1(n2245), .A2(n2436), .ZN(n2246) );
  AND3_X1 U2896 ( .A1(n4678), .A2(n2237), .A3(n2312), .ZN(n2247) );
  NOR2_X1 U2897 ( .A1(n4606), .A2(n4605), .ZN(n2248) );
  AND2_X1 U2898 ( .A1(n4066), .A2(n3638), .ZN(n2249) );
  NOR2_X1 U2899 ( .A1(n2745), .A2(n2427), .ZN(n2250) );
  NOR2_X1 U2900 ( .A1(n4064), .A2(n3790), .ZN(n2251) );
  NOR2_X1 U2901 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2252)
         );
  OR2_X1 U2902 ( .A1(n3819), .A2(n2402), .ZN(n2253) );
  NAND2_X1 U2903 ( .A1(n4067), .A2(n3861), .ZN(n2254) );
  INV_X1 U2904 ( .A(n3855), .ZN(n2413) );
  INV_X1 U2905 ( .A(IR_REG_28__SCAN_IN), .ZN(n2436) );
  INV_X1 U2906 ( .A(IR_REG_1__SCAN_IN), .ZN(n2362) );
  INV_X1 U2907 ( .A(IR_REG_0__SCAN_IN), .ZN(n2388) );
  INV_X1 U2908 ( .A(IR_REG_22__SCAN_IN), .ZN(n2487) );
  MUX2_X2 U2909 ( .A(n2512), .B(n2511), .S(n3095), .Z(n2552) );
  INV_X1 U2910 ( .A(n2357), .ZN(n2356) );
  NOR2_X1 U2911 ( .A1(n2358), .A2(n2360), .ZN(n2357) );
  NOR2_X1 U2912 ( .A1(n4058), .A2(n3888), .ZN(n2255) );
  AND2_X1 U2913 ( .A1(n2520), .A2(n2461), .ZN(n2522) );
  INV_X1 U2914 ( .A(n2320), .ZN(n4156) );
  NOR2_X1 U2915 ( .A1(n4233), .A2(n2321), .ZN(n2320) );
  NAND2_X1 U2916 ( .A1(n4212), .A2(n4424), .ZN(n2256) );
  XNOR2_X1 U2917 ( .A(n2935), .B(n2936), .ZN(n2257) );
  INV_X1 U2918 ( .A(n4271), .ZN(n2358) );
  AND2_X1 U2919 ( .A1(n2283), .A2(n2243), .ZN(n2520) );
  AND2_X1 U2920 ( .A1(n4185), .A2(n4170), .ZN(n2258) );
  NOR2_X1 U2921 ( .A1(n2244), .A2(n4260), .ZN(n2318) );
  INV_X1 U2922 ( .A(n2317), .ZN(n4313) );
  NOR2_X1 U2923 ( .A1(n4338), .A2(n4306), .ZN(n2317) );
  AND2_X1 U2924 ( .A1(n2313), .A2(n3518), .ZN(n2259) );
  AND2_X1 U2925 ( .A1(n3044), .A2(n2350), .ZN(n2260) );
  INV_X1 U2926 ( .A(n2372), .ZN(n2371) );
  NAND2_X1 U2927 ( .A1(n2241), .A2(n2448), .ZN(n2372) );
  AND2_X1 U2928 ( .A1(n2891), .A2(n2890), .ZN(n2261) );
  OR2_X1 U2929 ( .A1(n3053), .A2(n2258), .ZN(n2262) );
  INV_X1 U2930 ( .A(n3045), .ZN(n2361) );
  AND2_X1 U2931 ( .A1(n3223), .A2(n4708), .ZN(n2263) );
  INV_X1 U2932 ( .A(n3930), .ZN(n2301) );
  INV_X1 U2933 ( .A(n2424), .ZN(n2423) );
  NOR2_X1 U2934 ( .A1(n3868), .A2(n2257), .ZN(n2424) );
  OR2_X1 U2935 ( .A1(n2451), .A2(n2861), .ZN(n2264) );
  AND2_X1 U2936 ( .A1(n2936), .A2(n2935), .ZN(n2265) );
  NAND2_X1 U2937 ( .A1(n2421), .A2(n2952), .ZN(n2266) );
  OAI21_X1 U2938 ( .B1(n3415), .B2(n2251), .A(n3027), .ZN(n3532) );
  NAND2_X1 U2939 ( .A1(n2344), .A2(n2343), .ZN(n3357) );
  OAI21_X1 U2940 ( .B1(n3745), .B2(n2411), .A(n2410), .ZN(n3634) );
  NAND2_X1 U2941 ( .A1(n2346), .A2(n3023), .ZN(n3366) );
  OAI211_X1 U2942 ( .C1(n2393), .C2(n2971), .A(n2391), .B(n2389), .ZN(n2953)
         );
  INV_X1 U2943 ( .A(n4120), .ZN(n2336) );
  NAND2_X1 U2944 ( .A1(n2414), .A2(n2597), .ZN(n3776) );
  OR2_X1 U2945 ( .A1(n4713), .A2(REG1_REG_29__SCAN_IN), .ZN(n2267) );
  AND3_X1 U2946 ( .A1(n4678), .A2(n2237), .A3(n3339), .ZN(n2268) );
  NAND2_X1 U2947 ( .A1(n2552), .A2(DATAI_28_), .ZN(n4157) );
  INV_X1 U2948 ( .A(n4157), .ZN(n2324) );
  NAND2_X1 U2949 ( .A1(n2552), .A2(DATAI_26_), .ZN(n4199) );
  NAND2_X1 U2950 ( .A1(n2491), .A2(n2245), .ZN(n2989) );
  NAND2_X1 U2951 ( .A1(n2281), .A2(n2576), .ZN(n3249) );
  INV_X1 U2952 ( .A(IR_REG_24__SCAN_IN), .ZN(n2394) );
  AND2_X1 U2953 ( .A1(n3145), .A2(n4546), .ZN(n2269) );
  NAND2_X1 U2954 ( .A1(n2800), .A2(n2497), .ZN(n2270) );
  NAND2_X1 U2955 ( .A1(n2273), .A2(n2271), .ZN(n2528) );
  OR2_X1 U2956 ( .A1(n2800), .A2(n2761), .ZN(n2273) );
  NAND2_X1 U2957 ( .A1(n2274), .A2(n2663), .ZN(n3688) );
  AOI21_X2 U2958 ( .B1(n2277), .B2(n2276), .A(n2789), .ZN(n3759) );
  NOR2_X2 U2959 ( .A1(n2787), .A2(n2786), .ZN(n3878) );
  OAI21_X2 U2960 ( .B1(n2278), .B2(n2264), .A(n2862), .ZN(n3820) );
  NAND3_X1 U2961 ( .A1(n2388), .A2(n2279), .A3(n2362), .ZN(n2585) );
  NAND2_X2 U2962 ( .A1(n2506), .A2(n4539), .ZN(n2507) );
  NAND2_X1 U2963 ( .A1(n2282), .A2(n2698), .ZN(n3669) );
  NAND2_X1 U2964 ( .A1(n3787), .A2(n3788), .ZN(n2282) );
  INV_X1 U2965 ( .A(n2284), .ZN(n2887) );
  NAND2_X1 U2966 ( .A1(n4538), .A2(n3127), .ZN(n2284) );
  NAND2_X1 U2967 ( .A1(n2285), .A2(n2287), .ZN(n3076) );
  NAND2_X1 U2968 ( .A1(n4011), .A2(n2288), .ZN(n2285) );
  OR2_X1 U2969 ( .A1(n3088), .A2(n2294), .ZN(n2291) );
  NAND2_X1 U2970 ( .A1(n2291), .A2(n2292), .ZN(n4178) );
  NAND2_X2 U2971 ( .A1(n3932), .A2(n3935), .ZN(n3056) );
  NAND2_X1 U2972 ( .A1(n2468), .A2(IR_REG_31__SCAN_IN), .ZN(n2469) );
  OR2_X2 U2973 ( .A1(n3629), .A2(n2309), .ZN(n3111) );
  INV_X1 U2974 ( .A(n2318), .ZN(n4262) );
  AOI22_X1 U2975 ( .A1(n3209), .A2(n2328), .B1(n3145), .B2(n2327), .ZN(n2331)
         );
  INV_X1 U2976 ( .A(n2331), .ZN(n3178) );
  XNOR2_X2 U2977 ( .A(n2551), .B(IR_REG_1__SCAN_IN), .ZN(n4549) );
  NAND2_X1 U2978 ( .A1(n2387), .A2(IR_REG_31__SCAN_IN), .ZN(n2386) );
  NAND2_X1 U2979 ( .A1(n3337), .A2(n2337), .ZN(n2342) );
  NAND2_X1 U2980 ( .A1(n2342), .A2(n2341), .ZN(n3472) );
  NAND2_X1 U2981 ( .A1(n4345), .A2(n2348), .ZN(n2347) );
  INV_X1 U2982 ( .A(n2353), .ZN(n4243) );
  NOR2_X1 U2983 ( .A1(n2359), .A2(n2360), .ZN(n4269) );
  AND2_X1 U2984 ( .A1(n4308), .A2(n4440), .ZN(n2360) );
  NAND2_X1 U2985 ( .A1(n2388), .A2(n2362), .ZN(n2387) );
  NAND2_X1 U2986 ( .A1(n4193), .A2(n2368), .ZN(n2363) );
  NAND2_X1 U2987 ( .A1(n2363), .A2(n2365), .ZN(n3054) );
  AOI21_X1 U2988 ( .B1(n2373), .B2(n2448), .A(n3053), .ZN(n4169) );
  NOR2_X2 U2989 ( .A1(n2375), .A2(n2465), .ZN(n2374) );
  NAND2_X1 U2990 ( .A1(n2456), .A2(n2235), .ZN(n2375) );
  NAND2_X1 U2991 ( .A1(n3570), .A2(n2376), .ZN(n3037) );
  XNOR2_X2 U2992 ( .A(n2386), .B(IR_REG_2__SCAN_IN), .ZN(n4548) );
  NAND3_X1 U2993 ( .A1(n2409), .A2(n2407), .A3(n2411), .ZN(n2406) );
  NAND3_X1 U2994 ( .A1(n2414), .A2(n2597), .A3(n2611), .ZN(n3778) );
  AOI21_X1 U2995 ( .B1(n3870), .B2(n3867), .A(n3868), .ZN(n3644) );
  OAI211_X1 U2996 ( .C1(n3870), .C2(n2416), .A(n3883), .B(n2415), .ZN(n3014)
         );
  NAND2_X1 U2997 ( .A1(n3870), .A2(n2242), .ZN(n2415) );
  OAI21_X1 U2998 ( .B1(n2425), .B2(n2421), .A(n2418), .ZN(n2417) );
  INV_X1 U2999 ( .A(n2952), .ZN(n2425) );
  INV_X1 U3000 ( .A(n3834), .ZN(n3712) );
  NAND2_X1 U3001 ( .A1(n2753), .A2(n2431), .ZN(n2428) );
  INV_X1 U3002 ( .A(n2753), .ZN(n3810) );
  AND2_X1 U3003 ( .A1(n2491), .A2(n2466), .ZN(n2489) );
  INV_X1 U3004 ( .A(n2797), .ZN(n2438) );
  NAND2_X1 U3005 ( .A1(n2438), .A2(n2440), .ZN(n2488) );
  CLKBUF_X2 U3006 ( .A(n2557), .Z(n4070) );
  MUX2_X2 U3007 ( .A(REG0_REG_29__SCAN_IN), .B(n3111), .S(n4702), .Z(n3112) );
  NAND4_X1 U3008 ( .A1(n2584), .A2(n2583), .A3(n2582), .A4(n2581), .ZN(n2592)
         );
  NAND2_X1 U3009 ( .A1(n2598), .A2(REG1_REG_3__SCAN_IN), .ZN(n2583) );
  NAND2_X2 U3010 ( .A1(n3280), .A2(n4645), .ZN(n4648) );
  OAI211_X1 U3011 ( .C1(n3771), .C2(n2284), .A(n2889), .B(n2888), .ZN(n4212)
         );
  INV_X1 U3012 ( .A(n4350), .ZN(n3042) );
  INV_X1 U3013 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2790) );
  AND2_X1 U3014 ( .A1(n2836), .A2(n2835), .ZN(n2445) );
  OR2_X1 U3015 ( .A1(n4461), .A2(n3617), .ZN(n2446) );
  OR2_X1 U3016 ( .A1(n4288), .A2(n4276), .ZN(n2447) );
  NAND2_X1 U3017 ( .A1(n4409), .A2(n3872), .ZN(n2448) );
  OR2_X1 U3018 ( .A1(n4536), .A2(n4535), .ZN(U3499) );
  OR2_X1 U3019 ( .A1(n4473), .A2(n4472), .ZN(U3534) );
  OAI21_X1 U3020 ( .B1(n3759), .B2(n3755), .A(n3756), .ZN(n3845) );
  AND2_X1 U3021 ( .A1(n3702), .A2(n3703), .ZN(n2451) );
  OR2_X1 U3022 ( .A1(n4231), .A2(n4219), .ZN(n2452) );
  NAND2_X1 U3023 ( .A1(n2552), .A2(DATAI_24_), .ZN(n4424) );
  INV_X1 U3024 ( .A(n4424), .ZN(n4237) );
  OR2_X1 U3025 ( .A1(n3627), .A2(n4531), .ZN(n2453) );
  OR2_X1 U3026 ( .A1(n3627), .A2(n4467), .ZN(n2454) );
  OAI21_X1 U3027 ( .B1(n3688), .B2(n3689), .A(n3690), .ZN(n3787) );
  INV_X1 U3028 ( .A(IR_REG_4__SCAN_IN), .ZN(n2455) );
  NOR2_X1 U3029 ( .A1(n2485), .A2(IR_REG_19__SCAN_IN), .ZN(n2486) );
  OR2_X1 U3030 ( .A1(n2995), .A2(n4540), .ZN(n2981) );
  NAND2_X1 U3031 ( .A1(n4350), .A2(n3683), .ZN(n3043) );
  NAND2_X1 U3032 ( .A1(n3015), .A2(n3241), .ZN(n3935) );
  INV_X1 U3033 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2730) );
  AND2_X1 U3034 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n2476) );
  INV_X1 U3035 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4975) );
  OR2_X1 U3036 ( .A1(n2564), .A2(n2545), .ZN(n2550) );
  OR2_X1 U3037 ( .A1(n4350), .A2(n3683), .ZN(n3044) );
  INV_X1 U3038 ( .A(n4057), .ZN(n4461) );
  INV_X1 U3039 ( .A(n3837), .ZN(n3508) );
  INV_X1 U3040 ( .A(n3057), .ZN(n3320) );
  NOR2_X1 U3041 ( .A1(n2969), .A2(n3116), .ZN(n2496) );
  NAND2_X1 U3042 ( .A1(n2646), .A2(REG3_REG_7__SCAN_IN), .ZN(n2679) );
  OR2_X1 U3043 ( .A1(n2772), .A2(n5073), .ZN(n2791) );
  OR2_X1 U3044 ( .A1(n2791), .A2(n2790), .ZN(n2808) );
  OR2_X1 U3045 ( .A1(n2715), .A2(n3836), .ZN(n2731) );
  AND2_X1 U3046 ( .A1(n2634), .A2(REG3_REG_6__SCAN_IN), .ZN(n2646) );
  AND2_X1 U3047 ( .A1(n2998), .A2(n4645), .ZN(n3825) );
  AND2_X1 U3048 ( .A1(n2907), .A2(n2906), .ZN(n2925) );
  INV_X1 U3049 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3836) );
  INV_X1 U3050 ( .A(REG3_REG_16__SCAN_IN), .ZN(n5073) );
  OR2_X1 U3051 ( .A1(n2937), .A2(n4846), .ZN(n3626) );
  AND2_X1 U3052 ( .A1(n4179), .A2(n4157), .ZN(n3090) );
  NAND2_X1 U3053 ( .A1(n4273), .A2(n4296), .ZN(n3045) );
  AND2_X1 U3054 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2617) );
  OR2_X1 U3055 ( .A1(n3136), .A2(D_REG_0__SCAN_IN), .ZN(n2957) );
  INV_X1 U3056 ( .A(n4407), .ZN(n4170) );
  OR2_X1 U3057 ( .A1(n3136), .A2(n2968), .ZN(n3103) );
  OR3_X1 U3058 ( .A1(n2686), .A2(IR_REG_8__SCAN_IN), .A3(IR_REG_7__SCAN_IN), 
        .ZN(n2689) );
  INV_X1 U3059 ( .A(n4254), .ZN(n4260) );
  AND2_X1 U3060 ( .A1(n3010), .A2(n3009), .ZN(n3011) );
  AND2_X1 U3061 ( .A1(n2552), .A2(DATAI_21_), .ZN(n4296) );
  INV_X1 U3062 ( .A(n4199), .ZN(n3872) );
  OR2_X1 U3063 ( .A1(n2988), .A2(n2284), .ZN(n2944) );
  AND2_X1 U3064 ( .A1(n3147), .A2(n3146), .ZN(n4077) );
  AND2_X1 U3065 ( .A1(n4648), .A2(n4406), .ZN(n4382) );
  INV_X1 U3066 ( .A(n4385), .ZN(n4652) );
  INV_X1 U3067 ( .A(n4388), .ZN(n4196) );
  INV_X1 U3068 ( .A(n4645), .ZN(n4636) );
  NAND2_X1 U3069 ( .A1(n2957), .A2(n3139), .ZN(n3278) );
  INV_X1 U3070 ( .A(n4694), .ZN(n4474) );
  INV_X1 U3071 ( .A(n4468), .ZN(n4688) );
  INV_X1 U3072 ( .A(n3278), .ZN(n3109) );
  INV_X1 U3073 ( .A(n3275), .ZN(n3233) );
  AND2_X1 U3074 ( .A1(n2738), .A2(n2725), .ZN(n3443) );
  AND2_X1 U3075 ( .A1(n3147), .A2(n3135), .ZN(n4628) );
  AND2_X1 U3076 ( .A1(n3012), .A2(n3011), .ZN(n3013) );
  INV_X1 U3077 ( .A(n3883), .ZN(n3829) );
  NAND2_X1 U3078 ( .A1(n2944), .A2(n2943), .ZN(n4179) );
  NAND4_X1 U3079 ( .A1(n2828), .A2(n2827), .A3(n2826), .A4(n2825), .ZN(n4350)
         );
  NAND2_X1 U3080 ( .A1(n4077), .A2(n3189), .ZN(n4635) );
  NAND2_X1 U3081 ( .A1(n4648), .A2(n3359), .ZN(n4388) );
  AND2_X1 U3082 ( .A1(n3931), .A2(n3933), .ZN(n4671) );
  NAND2_X1 U3083 ( .A1(n4713), .A2(n4474), .ZN(n4467) );
  OR2_X1 U3084 ( .A1(n3110), .A2(n3278), .ZN(n4710) );
  NAND2_X1 U3085 ( .A1(n4702), .A2(n4474), .ZN(n4531) );
  AND3_X1 U3086 ( .A1(n4692), .A2(n4691), .A3(n4690), .ZN(n4709) );
  INV_X2 U3087 ( .A(n4700), .ZN(n4702) );
  NAND2_X1 U3088 ( .A1(n2495), .A2(n2494), .ZN(n3116) );
  INV_X1 U3089 ( .A(n3443), .ZN(n4667) );
  AND2_X1 U3090 ( .A1(n2625), .A2(n2624), .ZN(n4545) );
  NOR2_X1 U3091 ( .A1(n3114), .A2(n2536), .ZN(U4043) );
  NAND4_X1 U3092 ( .A1(n2484), .A2(n2464), .A3(n2463), .A4(n2462), .ZN(n2465)
         );
  NAND2_X1 U3093 ( .A1(n2991), .A2(n4797), .ZN(n2471) );
  NAND2_X2 U3094 ( .A1(n4538), .A2(n2478), .ZN(n2564) );
  NAND2_X1 U3095 ( .A1(n2598), .A2(REG1_REG_15__SCAN_IN), .ZN(n2483) );
  NAND2_X1 U3096 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2473) );
  NAND2_X1 U3097 ( .A1(n2699), .A2(REG3_REG_10__SCAN_IN), .ZN(n2715) );
  NAND2_X1 U3098 ( .A1(n2755), .A2(REG3_REG_14__SCAN_IN), .ZN(n2475) );
  INV_X1 U3099 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2474) );
  NAND2_X1 U3100 ( .A1(n2475), .A2(n2474), .ZN(n2477) );
  AND2_X1 U3101 ( .A1(n2477), .A2(n2772), .ZN(n3889) );
  NAND2_X1 U3102 ( .A1(n2600), .A2(n3889), .ZN(n2482) );
  NAND2_X1 U3103 ( .A1(n3895), .A2(REG0_REG_15__SCAN_IN), .ZN(n2481) );
  AND2_X1 U3104 ( .A1(n3127), .A2(n2479), .ZN(n2565) );
  NAND2_X1 U3105 ( .A1(n2840), .A2(REG2_REG_15__SCAN_IN), .ZN(n2480) );
  NAND4_X1 U3106 ( .A1(n2483), .A2(n2482), .A3(n2481), .A4(n2480), .ZN(n4058)
         );
  INV_X1 U3107 ( .A(n2484), .ZN(n2485) );
  OR2_X1 U3108 ( .A1(n2489), .A2(n2761), .ZN(n2490) );
  NOR2_X1 U3109 ( .A1(n2491), .A2(n2761), .ZN(n2492) );
  MUX2_X1 U3110 ( .A(n2761), .B(n2492), .S(IR_REG_25__SCAN_IN), .Z(n2493) );
  INV_X1 U3111 ( .A(n2489), .ZN(n2494) );
  XNOR2_X2 U3112 ( .A(n2499), .B(n2498), .ZN(n2506) );
  NAND2_X1 U3113 ( .A1(n2500), .A2(IR_REG_31__SCAN_IN), .ZN(n2501) );
  MUX2_X1 U3114 ( .A(IR_REG_31__SCAN_IN), .B(n2501), .S(IR_REG_21__SCAN_IN), 
        .Z(n2503) );
  INV_X1 U3115 ( .A(n2504), .ZN(n2502) );
  NAND2_X1 U3116 ( .A1(n2995), .A2(n2996), .ZN(n2975) );
  AND2_X2 U3117 ( .A1(n2553), .A2(n4694), .ZN(n2920) );
  NAND2_X1 U3118 ( .A1(n4058), .A2(n2920), .ZN(n2514) );
  BUF_X1 U3119 ( .A(n2770), .Z(n2933) );
  NAND2_X1 U3120 ( .A1(n2508), .A2(IR_REG_31__SCAN_IN), .ZN(n2509) );
  NAND2_X1 U3121 ( .A1(n2509), .A2(n4996), .ZN(n2778) );
  OR2_X1 U3122 ( .A1(n2509), .A2(n4996), .ZN(n2510) );
  NAND2_X1 U3123 ( .A1(n2436), .A2(n4799), .ZN(n2511) );
  MUX2_X1 U3124 ( .A(n4123), .B(DATAI_15_), .S(n3133), .Z(n3888) );
  NAND2_X1 U3125 ( .A1(n2913), .A2(n3888), .ZN(n2513) );
  NAND2_X1 U3126 ( .A1(n2514), .A2(n2513), .ZN(n3881) );
  NOR2_X1 U3127 ( .A1(n2733), .A2(REG3_REG_13__SCAN_IN), .ZN(n2515) );
  NOR2_X1 U3128 ( .A1(n2755), .A2(n2515), .ZN(n3814) );
  NAND2_X1 U3129 ( .A1(n2600), .A2(n3814), .ZN(n2519) );
  NAND2_X1 U3130 ( .A1(n2598), .A2(REG1_REG_13__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U3131 ( .A1(n2840), .A2(REG2_REG_13__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U3132 ( .A1(n3895), .A2(REG0_REG_13__SCAN_IN), .ZN(n2516) );
  NAND4_X1 U3133 ( .A1(n2519), .A2(n2518), .A3(n2517), .A4(n2516), .ZN(n4060)
         );
  NAND2_X1 U3134 ( .A1(n4060), .A2(n2913), .ZN(n2525) );
  NOR2_X1 U3135 ( .A1(n2520), .A2(n2761), .ZN(n2521) );
  MUX2_X1 U3136 ( .A(n2761), .B(n2521), .S(IR_REG_13__SCAN_IN), .Z(n2523) );
  OR2_X1 U3137 ( .A1(n2523), .A2(n2522), .ZN(n3440) );
  INV_X1 U3138 ( .A(n3440), .ZN(n4541) );
  MUX2_X1 U3139 ( .A(n4541), .B(DATAI_13_), .S(n3133), .Z(n3813) );
  NAND2_X1 U3140 ( .A1(n2899), .A2(n3813), .ZN(n2524) );
  NAND2_X1 U3141 ( .A1(n2525), .A2(n2524), .ZN(n2529) );
  OR2_X1 U3142 ( .A1(n2526), .A2(n4826), .ZN(n2527) );
  XNOR2_X1 U3143 ( .A(n2529), .B(n2233), .ZN(n3808) );
  NAND2_X1 U3144 ( .A1(n2887), .A2(REG3_REG_0__SCAN_IN), .ZN(n2532) );
  INV_X1 U3145 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2530) );
  AND2_X1 U3146 ( .A1(n2532), .A2(n2531), .ZN(n2534) );
  NAND2_X1 U3147 ( .A1(n2546), .A2(REG0_REG_0__SCAN_IN), .ZN(n2533) );
  NAND3_X2 U31480 ( .A1(n2535), .A2(n2534), .A3(n2533), .ZN(n4072) );
  NAND2_X1 U31490 ( .A1(n4072), .A2(n2984), .ZN(n2539) );
  MUX2_X1 U3150 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n3133), .Z(n3312) );
  NAND2_X1 U3151 ( .A1(n2553), .A2(n3312), .ZN(n2543) );
  INV_X1 U3152 ( .A(n2536), .ZN(n2540) );
  NAND2_X1 U3153 ( .A1(n2540), .A2(REG1_REG_0__SCAN_IN), .ZN(n2537) );
  AND2_X1 U3154 ( .A1(n2543), .A2(n2537), .ZN(n2538) );
  NAND2_X1 U3155 ( .A1(n2539), .A2(n2538), .ZN(n3187) );
  NAND2_X1 U3156 ( .A1(n4072), .A2(n2920), .ZN(n2542) );
  AOI22_X1 U3157 ( .A1(n2984), .A2(n3312), .B1(n2540), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2541) );
  NAND2_X1 U3158 ( .A1(n2542), .A2(n2541), .ZN(n3188) );
  NAND2_X1 U3159 ( .A1(n3187), .A2(n3188), .ZN(n3186) );
  NAND2_X1 U3160 ( .A1(n2543), .A2(n2917), .ZN(n2544) );
  NAND2_X1 U3161 ( .A1(n3186), .A2(n2544), .ZN(n3244) );
  INV_X1 U3162 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2545) );
  NAND2_X1 U3163 ( .A1(n2546), .A2(REG0_REG_1__SCAN_IN), .ZN(n2549) );
  NAND2_X1 U3164 ( .A1(n2565), .A2(REG2_REG_1__SCAN_IN), .ZN(n2548) );
  NAND2_X1 U3165 ( .A1(n2887), .A2(REG3_REG_1__SCAN_IN), .ZN(n2547) );
  NAND4_X1 U3166 ( .A1(n2550), .A2(n2549), .A3(n2548), .A4(n2547), .ZN(n2557)
         );
  NAND2_X1 U3167 ( .A1(n2557), .A2(n2984), .ZN(n2555) );
  NAND2_X1 U3168 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2551)
         );
  MUX2_X1 U3169 ( .A(n4549), .B(DATAI_1_), .S(n2552), .Z(n3241) );
  NAND2_X1 U3170 ( .A1(n2553), .A2(n3241), .ZN(n2554) );
  NAND2_X1 U3171 ( .A1(n2555), .A2(n2554), .ZN(n2556) );
  XNOR2_X1 U3172 ( .A(n2556), .B(n2233), .ZN(n2559) );
  NOR2_X1 U3173 ( .A1(n3286), .A2(n2770), .ZN(n2558) );
  AOI21_X1 U3174 ( .B1(n2557), .B2(n2920), .A(n2558), .ZN(n2560) );
  XNOR2_X1 U3175 ( .A(n2559), .B(n2560), .ZN(n3242) );
  NAND2_X1 U3176 ( .A1(n3244), .A2(n3242), .ZN(n3243) );
  INV_X1 U3177 ( .A(n2560), .ZN(n2561) );
  NAND2_X1 U3178 ( .A1(n2559), .A2(n2561), .ZN(n2562) );
  NAND2_X1 U3179 ( .A1(n3243), .A2(n2562), .ZN(n3251) );
  NAND2_X1 U3180 ( .A1(n2546), .A2(REG0_REG_2__SCAN_IN), .ZN(n2570) );
  INV_X1 U3181 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2563) );
  OR2_X1 U3182 ( .A1(n2564), .A2(n2563), .ZN(n2569) );
  NAND2_X1 U3183 ( .A1(n2565), .A2(REG2_REG_2__SCAN_IN), .ZN(n2567) );
  NAND2_X1 U3184 ( .A1(n2887), .A2(REG3_REG_2__SCAN_IN), .ZN(n2566) );
  AND2_X1 U3185 ( .A1(n2567), .A2(n2566), .ZN(n2568) );
  NAND2_X1 U3186 ( .A1(n2574), .A2(n2984), .ZN(n2572) );
  MUX2_X1 U3187 ( .A(n4548), .B(DATAI_2_), .S(n3133), .Z(n3106) );
  NAND2_X1 U3188 ( .A1(n2899), .A2(n3106), .ZN(n2571) );
  NAND2_X1 U3189 ( .A1(n2572), .A2(n2571), .ZN(n2573) );
  INV_X1 U3190 ( .A(n3106), .ZN(n3330) );
  NOR2_X1 U3191 ( .A1(n3330), .A2(n2770), .ZN(n2575) );
  AOI21_X1 U3192 ( .B1(n2574), .B2(n2920), .A(n2575), .ZN(n2577) );
  XNOR2_X1 U3193 ( .A(n2578), .B(n2577), .ZN(n3252) );
  INV_X1 U3194 ( .A(n3252), .ZN(n2576) );
  NAND2_X1 U3195 ( .A1(n2578), .A2(n2577), .ZN(n2579) );
  INV_X1 U3196 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2580) );
  NAND2_X1 U3197 ( .A1(n2600), .A2(n2580), .ZN(n2584) );
  NAND2_X1 U3198 ( .A1(n2840), .A2(REG2_REG_3__SCAN_IN), .ZN(n2582) );
  NAND2_X1 U3199 ( .A1(n2546), .A2(REG0_REG_3__SCAN_IN), .ZN(n2581) );
  NAND2_X1 U3200 ( .A1(n2592), .A2(n2984), .ZN(n2590) );
  NAND2_X1 U3201 ( .A1(n2585), .A2(IR_REG_31__SCAN_IN), .ZN(n2587) );
  NAND2_X1 U3202 ( .A1(n2587), .A2(n2586), .ZN(n2605) );
  OR2_X1 U3203 ( .A1(n2587), .A2(n2586), .ZN(n2588) );
  MUX2_X1 U3204 ( .A(n4547), .B(DATAI_3_), .S(n3133), .Z(n3262) );
  NAND2_X1 U3205 ( .A1(n2914), .A2(n3262), .ZN(n2589) );
  NAND2_X1 U3206 ( .A1(n2590), .A2(n2589), .ZN(n2591) );
  NOR2_X1 U3207 ( .A1(n3395), .A2(n2933), .ZN(n2593) );
  AOI21_X1 U3208 ( .B1(n2592), .B2(n2920), .A(n2593), .ZN(n2595) );
  XNOR2_X1 U3209 ( .A(n2594), .B(n2595), .ZN(n3258) );
  INV_X1 U32100 ( .A(n2594), .ZN(n2596) );
  NAND2_X1 U32110 ( .A1(n2596), .A2(n2595), .ZN(n2597) );
  NAND2_X1 U32120 ( .A1(n2598), .A2(REG1_REG_4__SCAN_IN), .ZN(n2604) );
  NOR2_X1 U32130 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2599) );
  NOR2_X1 U32140 ( .A1(n2617), .A2(n2599), .ZN(n3782) );
  NAND2_X1 U32150 ( .A1(n2600), .A2(n3782), .ZN(n2603) );
  NAND2_X1 U32160 ( .A1(n2546), .A2(REG0_REG_4__SCAN_IN), .ZN(n2602) );
  NAND2_X1 U32170 ( .A1(n2840), .A2(REG2_REG_4__SCAN_IN), .ZN(n2601) );
  NAND2_X1 U32180 ( .A1(n4069), .A2(n2984), .ZN(n2608) );
  NAND2_X1 U32190 ( .A1(n2605), .A2(IR_REG_31__SCAN_IN), .ZN(n2606) );
  XNOR2_X1 U32200 ( .A(n2606), .B(IR_REG_4__SCAN_IN), .ZN(n4546) );
  MUX2_X1 U32210 ( .A(n4546), .B(DATAI_4_), .S(n3133), .Z(n3781) );
  NAND2_X1 U32220 ( .A1(n2914), .A2(n3781), .ZN(n2607) );
  NAND2_X1 U32230 ( .A1(n2608), .A2(n2607), .ZN(n2609) );
  XNOR2_X1 U32240 ( .A(n2609), .B(n2917), .ZN(n2612) );
  INV_X1 U32250 ( .A(n3781), .ZN(n3297) );
  NOR2_X1 U32260 ( .A1(n3297), .A2(n2933), .ZN(n2610) );
  AOI21_X1 U32270 ( .B1(n4069), .B2(n2920), .A(n2610), .ZN(n2613) );
  XNOR2_X1 U32280 ( .A(n2612), .B(n2613), .ZN(n3777) );
  INV_X1 U32290 ( .A(n3777), .ZN(n2611) );
  INV_X1 U32300 ( .A(n2612), .ZN(n2615) );
  INV_X1 U32310 ( .A(n2613), .ZN(n2614) );
  NAND2_X1 U32320 ( .A1(n2615), .A2(n2614), .ZN(n2616) );
  NAND2_X1 U32330 ( .A1(n3778), .A2(n2616), .ZN(n3747) );
  NOR2_X1 U32340 ( .A1(n2617), .A2(REG3_REG_5__SCAN_IN), .ZN(n2618) );
  NOR2_X1 U32350 ( .A1(n2634), .A2(n2618), .ZN(n3750) );
  NAND2_X1 U32360 ( .A1(n2600), .A2(n3750), .ZN(n2622) );
  NAND2_X1 U32370 ( .A1(n2598), .A2(REG1_REG_5__SCAN_IN), .ZN(n2621) );
  NAND2_X1 U32380 ( .A1(n2840), .A2(REG2_REG_5__SCAN_IN), .ZN(n2620) );
  NAND2_X1 U32390 ( .A1(n2546), .A2(REG0_REG_5__SCAN_IN), .ZN(n2619) );
  NAND4_X1 U32400 ( .A1(n2622), .A2(n2621), .A3(n2620), .A4(n2619), .ZN(n4068)
         );
  NAND2_X1 U32410 ( .A1(n4068), .A2(n2913), .ZN(n2627) );
  NAND2_X1 U32420 ( .A1(n2375), .A2(IR_REG_31__SCAN_IN), .ZN(n2623) );
  MUX2_X1 U32430 ( .A(IR_REG_31__SCAN_IN), .B(n2623), .S(IR_REG_5__SCAN_IN), 
        .Z(n2625) );
  NOR2_X1 U32440 ( .A1(n2375), .A2(IR_REG_5__SCAN_IN), .ZN(n2653) );
  INV_X1 U32450 ( .A(n2653), .ZN(n2624) );
  MUX2_X1 U32460 ( .A(n4545), .B(DATAI_5_), .S(n3133), .Z(n3749) );
  NAND2_X1 U32470 ( .A1(n2899), .A2(n3749), .ZN(n2626) );
  NAND2_X1 U32480 ( .A1(n2627), .A2(n2626), .ZN(n2628) );
  XNOR2_X1 U32490 ( .A(n2628), .B(n2233), .ZN(n2632) );
  INV_X1 U32500 ( .A(n3749), .ZN(n3339) );
  NOR2_X1 U32510 ( .A1(n3339), .A2(n2933), .ZN(n2629) );
  AOI21_X1 U32520 ( .B1(n4068), .B2(n2920), .A(n2629), .ZN(n2630) );
  XNOR2_X1 U32530 ( .A(n2632), .B(n2630), .ZN(n3746) );
  INV_X1 U32540 ( .A(n2630), .ZN(n2631) );
  NAND2_X1 U32550 ( .A1(n2632), .A2(n2631), .ZN(n2633) );
  NAND2_X1 U32560 ( .A1(n2598), .A2(REG1_REG_6__SCAN_IN), .ZN(n2639) );
  NOR2_X1 U32570 ( .A1(n2634), .A2(REG3_REG_6__SCAN_IN), .ZN(n2635) );
  NOR2_X1 U32580 ( .A1(n2646), .A2(n2635), .ZN(n3862) );
  NAND2_X1 U32590 ( .A1(n2600), .A2(n3862), .ZN(n2638) );
  NAND2_X1 U32600 ( .A1(n2546), .A2(REG0_REG_6__SCAN_IN), .ZN(n2637) );
  NAND2_X1 U32610 ( .A1(n2840), .A2(REG2_REG_6__SCAN_IN), .ZN(n2636) );
  NAND4_X1 U32620 ( .A1(n2639), .A2(n2638), .A3(n2637), .A4(n2636), .ZN(n4067)
         );
  NAND2_X1 U32630 ( .A1(n4067), .A2(n2920), .ZN(n2642) );
  OR2_X1 U32640 ( .A1(n2653), .A2(n2761), .ZN(n2640) );
  XNOR2_X1 U32650 ( .A(n2640), .B(IR_REG_6__SCAN_IN), .ZN(n4544) );
  MUX2_X1 U32660 ( .A(n4544), .B(DATAI_6_), .S(n3133), .Z(n3861) );
  NAND2_X1 U32670 ( .A1(n2913), .A2(n3861), .ZN(n2641) );
  NAND2_X1 U32680 ( .A1(n2642), .A2(n2641), .ZN(n3855) );
  NAND2_X1 U32690 ( .A1(n4067), .A2(n2984), .ZN(n2644) );
  NAND2_X1 U32700 ( .A1(n2899), .A2(n3861), .ZN(n2643) );
  NAND2_X1 U32710 ( .A1(n2644), .A2(n2643), .ZN(n2645) );
  XNOR2_X1 U32720 ( .A(n2645), .B(n2234), .ZN(n3856) );
  NAND2_X1 U32730 ( .A1(n2598), .A2(REG1_REG_7__SCAN_IN), .ZN(n2652) );
  INV_X1 U32740 ( .A(n2646), .ZN(n2647) );
  INV_X1 U32750 ( .A(REG3_REG_7__SCAN_IN), .ZN(n3221) );
  NAND2_X1 U32760 ( .A1(n2647), .A2(n3221), .ZN(n2648) );
  AND2_X1 U32770 ( .A1(n2648), .A2(n2679), .ZN(n3639) );
  NAND2_X1 U32780 ( .A1(n2600), .A2(n3639), .ZN(n2651) );
  NAND2_X1 U32790 ( .A1(n2546), .A2(REG0_REG_7__SCAN_IN), .ZN(n2650) );
  NAND2_X1 U32800 ( .A1(n2840), .A2(REG2_REG_7__SCAN_IN), .ZN(n2649) );
  NAND4_X1 U32810 ( .A1(n2652), .A2(n2651), .A3(n2650), .A4(n2649), .ZN(n4066)
         );
  NAND2_X1 U32820 ( .A1(n4066), .A2(n2913), .ZN(n2657) );
  NAND2_X1 U32830 ( .A1(n2653), .A2(n5011), .ZN(n2686) );
  NAND2_X1 U32840 ( .A1(n2686), .A2(IR_REG_31__SCAN_IN), .ZN(n2654) );
  NAND2_X1 U32850 ( .A1(n2654), .A2(n4798), .ZN(n2668) );
  OR2_X1 U32860 ( .A1(n2654), .A2(n4798), .ZN(n2655) );
  MUX2_X1 U32870 ( .A(n4543), .B(DATAI_7_), .S(n3133), .Z(n3638) );
  NAND2_X1 U32880 ( .A1(n2914), .A2(n3638), .ZN(n2656) );
  NAND2_X1 U32890 ( .A1(n2657), .A2(n2656), .ZN(n2658) );
  XNOR2_X1 U32900 ( .A(n2658), .B(n2233), .ZN(n2662) );
  NOR2_X1 U32910 ( .A1(n3360), .A2(n2933), .ZN(n2659) );
  AOI21_X1 U32920 ( .B1(n4066), .B2(n2920), .A(n2659), .ZN(n2660) );
  XNOR2_X1 U32930 ( .A(n2662), .B(n2660), .ZN(n3635) );
  INV_X1 U32940 ( .A(n2660), .ZN(n2661) );
  NAND2_X1 U32950 ( .A1(n2662), .A2(n2661), .ZN(n2663) );
  XNOR2_X1 U32960 ( .A(n2679), .B(REG3_REG_8__SCAN_IN), .ZN(n4644) );
  NAND2_X1 U32970 ( .A1(n2600), .A2(n4644), .ZN(n2667) );
  NAND2_X1 U32980 ( .A1(n2598), .A2(REG1_REG_8__SCAN_IN), .ZN(n2666) );
  NAND2_X1 U32990 ( .A1(n2840), .A2(REG2_REG_8__SCAN_IN), .ZN(n2665) );
  NAND2_X1 U33000 ( .A1(n3895), .A2(REG0_REG_8__SCAN_IN), .ZN(n2664) );
  NAND4_X1 U33010 ( .A1(n2667), .A2(n2666), .A3(n2665), .A4(n2664), .ZN(n4065)
         );
  NAND2_X1 U33020 ( .A1(n4065), .A2(n2913), .ZN(n2671) );
  NAND2_X1 U33030 ( .A1(n2668), .A2(IR_REG_31__SCAN_IN), .ZN(n2669) );
  XNOR2_X1 U33040 ( .A(n2669), .B(IR_REG_8__SCAN_IN), .ZN(n4542) );
  MUX2_X1 U33050 ( .A(n4542), .B(DATAI_8_), .S(n3133), .Z(n3696) );
  NAND2_X1 U33060 ( .A1(n2899), .A2(n3696), .ZN(n2670) );
  NAND2_X1 U33070 ( .A1(n2671), .A2(n2670), .ZN(n2672) );
  XNOR2_X1 U33080 ( .A(n2672), .B(n2234), .ZN(n2675) );
  NAND2_X1 U33090 ( .A1(n4065), .A2(n2920), .ZN(n2674) );
  NAND2_X1 U33100 ( .A1(n2984), .A2(n3696), .ZN(n2673) );
  NAND2_X1 U33110 ( .A1(n2674), .A2(n2673), .ZN(n2676) );
  AND2_X1 U33120 ( .A1(n2675), .A2(n2676), .ZN(n3689) );
  INV_X1 U33130 ( .A(n2675), .ZN(n2678) );
  INV_X1 U33140 ( .A(n2676), .ZN(n2677) );
  NAND2_X1 U33150 ( .A1(n2678), .A2(n2677), .ZN(n3690) );
  INV_X1 U33160 ( .A(n2679), .ZN(n2680) );
  AOI21_X1 U33170 ( .B1(n2680), .B2(REG3_REG_8__SCAN_IN), .A(
        REG3_REG_9__SCAN_IN), .ZN(n2681) );
  OR2_X1 U33180 ( .A1(n2681), .A2(n2699), .ZN(n3418) );
  INV_X1 U33190 ( .A(n3418), .ZN(n3791) );
  NAND2_X1 U33200 ( .A1(n2600), .A2(n3791), .ZN(n2685) );
  NAND2_X1 U33210 ( .A1(n2598), .A2(REG1_REG_9__SCAN_IN), .ZN(n2684) );
  NAND2_X1 U33220 ( .A1(n3895), .A2(REG0_REG_9__SCAN_IN), .ZN(n2683) );
  NAND2_X1 U33230 ( .A1(n2840), .A2(REG2_REG_9__SCAN_IN), .ZN(n2682) );
  NAND4_X1 U33240 ( .A1(n2685), .A2(n2684), .A3(n2683), .A4(n2682), .ZN(n4064)
         );
  NAND2_X1 U33250 ( .A1(n4064), .A2(n2913), .ZN(n2692) );
  NAND2_X1 U33260 ( .A1(n2689), .A2(IR_REG_31__SCAN_IN), .ZN(n2687) );
  MUX2_X1 U33270 ( .A(IR_REG_31__SCAN_IN), .B(n2687), .S(IR_REG_9__SCAN_IN), 
        .Z(n2688) );
  INV_X1 U33280 ( .A(n2688), .ZN(n2690) );
  MUX2_X1 U33290 ( .A(n4553), .B(DATAI_9_), .S(n3133), .Z(n3790) );
  NAND2_X1 U33300 ( .A1(n2914), .A2(n3790), .ZN(n2691) );
  NAND2_X1 U33310 ( .A1(n2692), .A2(n2691), .ZN(n2693) );
  XNOR2_X1 U33320 ( .A(n2693), .B(n2233), .ZN(n2695) );
  INV_X1 U33330 ( .A(n3790), .ZN(n3459) );
  NOR2_X1 U33340 ( .A1(n3459), .A2(n2946), .ZN(n2694) );
  AOI21_X1 U33350 ( .B1(n4064), .B2(n2920), .A(n2694), .ZN(n2696) );
  XNOR2_X1 U33360 ( .A(n2695), .B(n2696), .ZN(n3788) );
  INV_X1 U33370 ( .A(n2695), .ZN(n2697) );
  NAND2_X1 U33380 ( .A1(n2697), .A2(n2696), .ZN(n2698) );
  OR2_X1 U33390 ( .A1(n2699), .A2(REG3_REG_10__SCAN_IN), .ZN(n2700) );
  AND2_X1 U33400 ( .A1(n2715), .A2(n2700), .ZN(n4637) );
  NAND2_X1 U33410 ( .A1(n2600), .A2(n4637), .ZN(n2704) );
  NAND2_X1 U33420 ( .A1(n2598), .A2(REG1_REG_10__SCAN_IN), .ZN(n2703) );
  NAND2_X1 U33430 ( .A1(n3895), .A2(REG0_REG_10__SCAN_IN), .ZN(n2702) );
  NAND2_X1 U33440 ( .A1(n2840), .A2(REG2_REG_10__SCAN_IN), .ZN(n2701) );
  NAND4_X1 U33450 ( .A1(n2704), .A2(n2703), .A3(n2702), .A4(n2701), .ZN(n4063)
         );
  NAND2_X1 U33460 ( .A1(n4063), .A2(n2913), .ZN(n2707) );
  OR2_X1 U33470 ( .A1(n2721), .A2(n2761), .ZN(n2705) );
  XNOR2_X1 U33480 ( .A(n2705), .B(IR_REG_10__SCAN_IN), .ZN(n3448) );
  MUX2_X1 U33490 ( .A(n3448), .B(DATAI_10_), .S(n3133), .Z(n3674) );
  NAND2_X1 U33500 ( .A1(n2899), .A2(n3674), .ZN(n2706) );
  NAND2_X1 U33510 ( .A1(n2707), .A2(n2706), .ZN(n2708) );
  XNOR2_X1 U33520 ( .A(n2708), .B(n2917), .ZN(n2710) );
  NOR2_X1 U3353 ( .A1(n3534), .A2(n2946), .ZN(n2709) );
  AOI21_X1 U33540 ( .B1(n4063), .B2(n2920), .A(n2709), .ZN(n2711) );
  XNOR2_X1 U3355 ( .A(n2710), .B(n2711), .ZN(n3670) );
  INV_X1 U3356 ( .A(n2710), .ZN(n2713) );
  INV_X1 U3357 ( .A(n2711), .ZN(n2712) );
  NAND2_X1 U3358 ( .A1(n2713), .A2(n2712), .ZN(n2714) );
  NAND2_X1 U3359 ( .A1(n2715), .A2(n3836), .ZN(n2716) );
  AND2_X1 U3360 ( .A1(n2731), .A2(n2716), .ZN(n3838) );
  NAND2_X1 U3361 ( .A1(n2600), .A2(n3838), .ZN(n2720) );
  NAND2_X1 U3362 ( .A1(n2598), .A2(REG1_REG_11__SCAN_IN), .ZN(n2719) );
  NAND2_X1 U3363 ( .A1(n2840), .A2(REG2_REG_11__SCAN_IN), .ZN(n2718) );
  NAND2_X1 U3364 ( .A1(n3895), .A2(REG0_REG_11__SCAN_IN), .ZN(n2717) );
  NAND4_X1 U3365 ( .A1(n2720), .A2(n2719), .A3(n2718), .A4(n2717), .ZN(n4062)
         );
  NAND2_X1 U3366 ( .A1(n4062), .A2(n2913), .ZN(n2727) );
  NAND2_X1 U3367 ( .A1(n2721), .A2(n5001), .ZN(n2722) );
  NAND2_X1 U3368 ( .A1(n2722), .A2(IR_REG_31__SCAN_IN), .ZN(n2724) );
  INV_X1 U3369 ( .A(IR_REG_11__SCAN_IN), .ZN(n2723) );
  NAND2_X1 U3370 ( .A1(n2724), .A2(n2723), .ZN(n2738) );
  OR2_X1 U3371 ( .A1(n2724), .A2(n2723), .ZN(n2725) );
  MUX2_X1 U3372 ( .A(n3443), .B(DATAI_11_), .S(n3133), .Z(n3837) );
  NAND2_X1 U3373 ( .A1(n2899), .A2(n3837), .ZN(n2726) );
  NAND2_X1 U3374 ( .A1(n2727), .A2(n2726), .ZN(n2728) );
  XNOR2_X1 U3375 ( .A(n2728), .B(n2917), .ZN(n3832) );
  NOR2_X1 U3376 ( .A1(n3508), .A2(n2946), .ZN(n2729) );
  AOI21_X1 U3377 ( .B1(n4062), .B2(n2920), .A(n2729), .ZN(n3831) );
  NAND2_X1 U3378 ( .A1(n2598), .A2(REG1_REG_12__SCAN_IN), .ZN(n2737) );
  AND2_X1 U3379 ( .A1(n2731), .A2(n2730), .ZN(n2732) );
  NOR2_X1 U3380 ( .A1(n2733), .A2(n2732), .ZN(n3721) );
  NAND2_X1 U3381 ( .A1(n2600), .A2(n3721), .ZN(n2736) );
  NAND2_X1 U3382 ( .A1(n3895), .A2(REG0_REG_12__SCAN_IN), .ZN(n2735) );
  NAND2_X1 U3383 ( .A1(n2840), .A2(REG2_REG_12__SCAN_IN), .ZN(n2734) );
  NAND4_X1 U3384 ( .A1(n2737), .A2(n2736), .A3(n2735), .A4(n2734), .ZN(n4061)
         );
  NAND2_X1 U3385 ( .A1(n4061), .A2(n2913), .ZN(n2741) );
  NAND2_X1 U3386 ( .A1(n2738), .A2(IR_REG_31__SCAN_IN), .ZN(n2739) );
  XNOR2_X1 U3387 ( .A(n2739), .B(IR_REG_12__SCAN_IN), .ZN(n3452) );
  MUX2_X1 U3388 ( .A(n3452), .B(DATAI_12_), .S(n3133), .Z(n3720) );
  NAND2_X1 U3389 ( .A1(n2914), .A2(n3720), .ZN(n2740) );
  NAND2_X1 U3390 ( .A1(n2741), .A2(n2740), .ZN(n2742) );
  XNOR2_X1 U3391 ( .A(n2742), .B(n2234), .ZN(n2746) );
  NAND2_X1 U3392 ( .A1(n4061), .A2(n2920), .ZN(n2744) );
  NAND2_X1 U3393 ( .A1(n2913), .A2(n3720), .ZN(n2743) );
  NAND2_X1 U3394 ( .A1(n2744), .A2(n2743), .ZN(n2747) );
  NAND2_X1 U3395 ( .A1(n2746), .A2(n2747), .ZN(n3715) );
  OAI21_X1 U3396 ( .B1(n3832), .B2(n3831), .A(n3715), .ZN(n2745) );
  NAND3_X1 U3397 ( .A1(n3715), .A2(n3831), .A3(n3832), .ZN(n2750) );
  INV_X1 U3398 ( .A(n2746), .ZN(n2749) );
  INV_X1 U3399 ( .A(n2747), .ZN(n2748) );
  NAND2_X1 U3400 ( .A1(n2749), .A2(n2748), .ZN(n3714) );
  AND2_X1 U3401 ( .A1(n2750), .A2(n3714), .ZN(n2751) );
  INV_X1 U3402 ( .A(n4060), .ZN(n3577) );
  INV_X1 U3403 ( .A(n3813), .ZN(n3518) );
  OAI22_X1 U3404 ( .A1(n3577), .A2(n2947), .B1(n2946), .B2(n3518), .ZN(n3807)
         );
  INV_X1 U3405 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2754) );
  XNOR2_X1 U3406 ( .A(n2755), .B(n2754), .ZN(n3657) );
  NAND2_X1 U3407 ( .A1(n2600), .A2(n3657), .ZN(n2759) );
  NAND2_X1 U3408 ( .A1(n2598), .A2(REG1_REG_14__SCAN_IN), .ZN(n2758) );
  NAND2_X1 U3409 ( .A1(n2840), .A2(REG2_REG_14__SCAN_IN), .ZN(n2757) );
  NAND2_X1 U3410 ( .A1(n3895), .A2(REG0_REG_14__SCAN_IN), .ZN(n2756) );
  NAND4_X1 U3411 ( .A1(n2759), .A2(n2758), .A3(n2757), .A4(n2756), .ZN(n4059)
         );
  NAND2_X1 U3412 ( .A1(n4059), .A2(n2913), .ZN(n2765) );
  NOR2_X1 U3413 ( .A1(n2522), .A2(n2761), .ZN(n2760) );
  MUX2_X1 U3414 ( .A(n2761), .B(n2760), .S(IR_REG_14__SCAN_IN), .Z(n2762) );
  INV_X1 U3415 ( .A(n2762), .ZN(n2763) );
  AND2_X1 U3416 ( .A1(n2508), .A2(n2763), .ZN(n4120) );
  MUX2_X1 U3417 ( .A(n4120), .B(DATAI_14_), .S(n3133), .Z(n3656) );
  NAND2_X1 U3418 ( .A1(n2899), .A2(n3656), .ZN(n2764) );
  NAND2_X1 U3419 ( .A1(n2765), .A2(n2764), .ZN(n2766) );
  XNOR2_X1 U3420 ( .A(n2766), .B(n2917), .ZN(n2769) );
  NOR2_X1 U3421 ( .A1(n3581), .A2(n2946), .ZN(n2767) );
  AOI21_X1 U3422 ( .B1(n4059), .B2(n2920), .A(n2767), .ZN(n2768) );
  NOR2_X1 U3423 ( .A1(n2769), .A2(n2768), .ZN(n3650) );
  NAND2_X1 U3424 ( .A1(n2769), .A2(n2768), .ZN(n3651) );
  INV_X1 U3425 ( .A(n4058), .ZN(n3073) );
  INV_X1 U3426 ( .A(n3888), .ZN(n3594) );
  OAI22_X1 U3427 ( .A1(n3073), .A2(n2770), .B1(n2945), .B2(n3594), .ZN(n2771)
         );
  XOR2_X1 U3428 ( .A(n2234), .B(n2771), .Z(n2786) );
  NAND2_X1 U3429 ( .A1(n2787), .A2(n2786), .ZN(n3879) );
  NAND2_X1 U3430 ( .A1(n2772), .A2(n5073), .ZN(n2773) );
  AND2_X1 U3431 ( .A1(n2791), .A2(n2773), .ZN(n3740) );
  NAND2_X1 U3432 ( .A1(n2600), .A2(n3740), .ZN(n2777) );
  NAND2_X1 U3433 ( .A1(n2598), .A2(REG1_REG_16__SCAN_IN), .ZN(n2776) );
  NAND2_X1 U3434 ( .A1(n2840), .A2(REG2_REG_16__SCAN_IN), .ZN(n2775) );
  NAND2_X1 U3435 ( .A1(n3895), .A2(REG0_REG_16__SCAN_IN), .ZN(n2774) );
  NAND4_X1 U3436 ( .A1(n2777), .A2(n2776), .A3(n2775), .A4(n2774), .ZN(n4057)
         );
  NAND2_X1 U3437 ( .A1(n4057), .A2(n2913), .ZN(n2781) );
  NAND2_X1 U3438 ( .A1(n2778), .A2(IR_REG_31__SCAN_IN), .ZN(n2779) );
  XNOR2_X1 U3439 ( .A(n2779), .B(IR_REG_16__SCAN_IN), .ZN(n4124) );
  MUX2_X1 U3440 ( .A(n4124), .B(DATAI_16_), .S(n3133), .Z(n3739) );
  NAND2_X1 U3441 ( .A1(n2914), .A2(n3739), .ZN(n2780) );
  NAND2_X1 U3442 ( .A1(n2781), .A2(n2780), .ZN(n2782) );
  XNOR2_X1 U3443 ( .A(n2782), .B(n2917), .ZN(n2785) );
  INV_X1 U3444 ( .A(n3739), .ZN(n3617) );
  NOR2_X1 U3445 ( .A1(n3617), .A2(n2946), .ZN(n2783) );
  AOI21_X1 U3446 ( .B1(n4057), .B2(n2920), .A(n2783), .ZN(n2784) );
  NAND2_X1 U3447 ( .A1(n2785), .A2(n2784), .ZN(n2788) );
  OAI21_X1 U3448 ( .B1(n2785), .B2(n2784), .A(n2788), .ZN(n3737) );
  INV_X1 U3449 ( .A(n2788), .ZN(n2789) );
  NAND2_X1 U3450 ( .A1(n2598), .A2(REG1_REG_17__SCAN_IN), .ZN(n2796) );
  NAND2_X1 U3451 ( .A1(n2791), .A2(n2790), .ZN(n2792) );
  AND2_X1 U3452 ( .A1(n2808), .A2(n2792), .ZN(n4377) );
  NAND2_X1 U3453 ( .A1(n2600), .A2(n4377), .ZN(n2795) );
  NAND2_X1 U3454 ( .A1(n3895), .A2(REG0_REG_17__SCAN_IN), .ZN(n2794) );
  NAND2_X1 U3455 ( .A1(n2840), .A2(REG2_REG_17__SCAN_IN), .ZN(n2793) );
  NAND4_X1 U3456 ( .A1(n2796), .A2(n2795), .A3(n2794), .A4(n2793), .ZN(n4056)
         );
  NAND2_X1 U3457 ( .A1(n4056), .A2(n2913), .ZN(n2803) );
  NAND2_X1 U34580 ( .A1(n2797), .A2(IR_REG_31__SCAN_IN), .ZN(n2798) );
  MUX2_X1 U34590 ( .A(IR_REG_31__SCAN_IN), .B(n2798), .S(IR_REG_17__SCAN_IN), 
        .Z(n2799) );
  INV_X1 U3460 ( .A(n2799), .ZN(n2801) );
  NOR2_X1 U3461 ( .A1(n2801), .A2(n2800), .ZN(n4127) );
  INV_X1 U3462 ( .A(n4127), .ZN(n4662) );
  INV_X1 U3463 ( .A(DATAI_17_), .ZN(n4661) );
  MUX2_X1 U3464 ( .A(n4662), .B(n4661), .S(n3133), .Z(n4458) );
  NAND2_X1 U3465 ( .A1(n2914), .A2(n4383), .ZN(n2802) );
  NAND2_X1 U3466 ( .A1(n2803), .A2(n2802), .ZN(n2804) );
  XNOR2_X1 U34670 ( .A(n2804), .B(n2917), .ZN(n2807) );
  NOR2_X1 U3468 ( .A1(n2946), .A2(n4458), .ZN(n2805) );
  AOI21_X1 U34690 ( .B1(n4056), .B2(n2920), .A(n2805), .ZN(n2806) );
  NOR2_X1 U3470 ( .A1(n2807), .A2(n2806), .ZN(n3755) );
  NAND2_X1 U34710 ( .A1(n2807), .A2(n2806), .ZN(n3756) );
  NAND2_X1 U3472 ( .A1(n2598), .A2(REG1_REG_18__SCAN_IN), .ZN(n2813) );
  AND2_X1 U34730 ( .A1(n2808), .A2(n3850), .ZN(n2809) );
  NOR2_X1 U3474 ( .A1(n2838), .A2(n2809), .ZN(n4358) );
  NAND2_X1 U34750 ( .A1(n2600), .A2(n4358), .ZN(n2812) );
  NAND2_X1 U3476 ( .A1(n3895), .A2(REG0_REG_18__SCAN_IN), .ZN(n2811) );
  NAND2_X1 U34770 ( .A1(n2840), .A2(REG2_REG_18__SCAN_IN), .ZN(n2810) );
  NAND4_X1 U3478 ( .A1(n2813), .A2(n2812), .A3(n2811), .A4(n2810), .ZN(n4370)
         );
  NAND2_X1 U34790 ( .A1(n4370), .A2(n2913), .ZN(n2817) );
  INV_X1 U3480 ( .A(n2800), .ZN(n2814) );
  NAND2_X1 U34810 ( .A1(n2814), .A2(IR_REG_31__SCAN_IN), .ZN(n2815) );
  MUX2_X1 U3482 ( .A(n4138), .B(DATAI_18_), .S(n3133), .Z(n4349) );
  NAND2_X1 U34830 ( .A1(n2899), .A2(n4349), .ZN(n2816) );
  NAND2_X1 U3484 ( .A1(n2817), .A2(n2816), .ZN(n2818) );
  XNOR2_X1 U34850 ( .A(n2818), .B(n2234), .ZN(n2821) );
  NAND2_X1 U3486 ( .A1(n4370), .A2(n2920), .ZN(n2820) );
  NAND2_X1 U34870 ( .A1(n2913), .A2(n4349), .ZN(n2819) );
  NAND2_X1 U3488 ( .A1(n2820), .A2(n2819), .ZN(n2822) );
  NAND2_X1 U34890 ( .A1(n2821), .A2(n2822), .ZN(n3847) );
  NAND2_X1 U3490 ( .A1(n3845), .A2(n3847), .ZN(n3844) );
  INV_X1 U34910 ( .A(n2821), .ZN(n2824) );
  INV_X1 U3492 ( .A(n2822), .ZN(n2823) );
  NAND2_X1 U34930 ( .A1(n2824), .A2(n2823), .ZN(n3846) );
  NAND2_X1 U3494 ( .A1(n3844), .A2(n3846), .ZN(n3680) );
  INV_X1 U34950 ( .A(REG3_REG_19__SCAN_IN), .ZN(n5069) );
  XNOR2_X1 U3496 ( .A(n2838), .B(n5069), .ZN(n4339) );
  NAND2_X1 U34970 ( .A1(n2600), .A2(n4339), .ZN(n2828) );
  NAND2_X1 U3498 ( .A1(n2598), .A2(REG1_REG_19__SCAN_IN), .ZN(n2827) );
  NAND2_X1 U34990 ( .A1(n2840), .A2(REG2_REG_19__SCAN_IN), .ZN(n2826) );
  NAND2_X1 U3500 ( .A1(n3895), .A2(REG0_REG_19__SCAN_IN), .ZN(n2825) );
  INV_X1 U35010 ( .A(DATAI_19_), .ZN(n2829) );
  MUX2_X1 U3502 ( .A(n4144), .B(n2829), .S(n2552), .Z(n4336) );
  OAI22_X1 U35030 ( .A1(n3042), .A2(n2947), .B1(n2946), .B2(n4336), .ZN(n2834)
         );
  NAND2_X1 U3504 ( .A1(n4350), .A2(n2913), .ZN(n2831) );
  INV_X1 U35050 ( .A(n4336), .ZN(n3683) );
  NAND2_X1 U35060 ( .A1(n2914), .A2(n3683), .ZN(n2830) );
  NAND2_X1 U35070 ( .A1(n2831), .A2(n2830), .ZN(n2832) );
  XNOR2_X1 U35080 ( .A(n2832), .B(n2233), .ZN(n2833) );
  XOR2_X1 U35090 ( .A(n2834), .B(n2833), .Z(n3679) );
  INV_X1 U35100 ( .A(n2833), .ZN(n2836) );
  INV_X1 U35110 ( .A(n2834), .ZN(n2835) );
  AOI21_X1 U35120 ( .B1(n3680), .B2(n3679), .A(n2445), .ZN(n3701) );
  AND2_X1 U35130 ( .A1(REG3_REG_19__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2837) );
  AOI21_X1 U35140 ( .B1(n2838), .B2(REG3_REG_19__SCAN_IN), .A(
        REG3_REG_20__SCAN_IN), .ZN(n2839) );
  OR2_X1 U35150 ( .A1(n2849), .A2(n2839), .ZN(n4316) );
  INV_X1 U35160 ( .A(n4316), .ZN(n3802) );
  NAND2_X1 U35170 ( .A1(n2600), .A2(n3802), .ZN(n2844) );
  NAND2_X1 U35180 ( .A1(n2598), .A2(REG1_REG_20__SCAN_IN), .ZN(n2843) );
  NAND2_X1 U35190 ( .A1(n3895), .A2(REG0_REG_20__SCAN_IN), .ZN(n2842) );
  NAND2_X1 U35200 ( .A1(n2840), .A2(REG2_REG_20__SCAN_IN), .ZN(n2841) );
  NAND4_X1 U35210 ( .A1(n2844), .A2(n2843), .A3(n2842), .A4(n2841), .ZN(n4055)
         );
  NAND2_X1 U35220 ( .A1(n4055), .A2(n2913), .ZN(n2846) );
  NAND2_X1 U35230 ( .A1(n2914), .A2(n4306), .ZN(n2845) );
  NAND2_X1 U35240 ( .A1(n2846), .A2(n2845), .ZN(n2847) );
  XNOR2_X1 U35250 ( .A(n2847), .B(n2917), .ZN(n2860) );
  INV_X1 U35260 ( .A(n4306), .ZN(n4314) );
  NOR2_X1 U35270 ( .A1(n2946), .A2(n4314), .ZN(n2848) );
  AOI21_X1 U35280 ( .B1(n4055), .B2(n2920), .A(n2848), .ZN(n2859) );
  NOR2_X1 U35290 ( .A1(n2860), .A2(n2859), .ZN(n3796) );
  OR2_X1 U35300 ( .A1(n2849), .A2(REG3_REG_21__SCAN_IN), .ZN(n2850) );
  AND2_X1 U35310 ( .A1(n2850), .A2(n2873), .ZN(n4293) );
  NAND2_X1 U35320 ( .A1(n2600), .A2(n4293), .ZN(n2854) );
  NAND2_X1 U35330 ( .A1(n2598), .A2(REG1_REG_21__SCAN_IN), .ZN(n2853) );
  NAND2_X1 U35340 ( .A1(n2840), .A2(REG2_REG_21__SCAN_IN), .ZN(n2852) );
  NAND2_X1 U35350 ( .A1(n3895), .A2(REG0_REG_21__SCAN_IN), .ZN(n2851) );
  NAND4_X1 U35360 ( .A1(n2854), .A2(n2853), .A3(n2852), .A4(n2851), .ZN(n4273)
         );
  NAND2_X1 U35370 ( .A1(n4273), .A2(n2913), .ZN(n2856) );
  NAND2_X1 U35380 ( .A1(n2914), .A2(n4296), .ZN(n2855) );
  NAND2_X1 U35390 ( .A1(n2856), .A2(n2855), .ZN(n2857) );
  XNOR2_X1 U35400 ( .A(n2857), .B(n2917), .ZN(n3702) );
  NOR2_X1 U35410 ( .A1(n2946), .A2(n4440), .ZN(n2858) );
  AOI21_X1 U35420 ( .B1(n4273), .B2(n2920), .A(n2858), .ZN(n3703) );
  NAND2_X1 U35430 ( .A1(n2860), .A2(n2859), .ZN(n3797) );
  XNOR2_X1 U35440 ( .A(n2873), .B(REG3_REG_22__SCAN_IN), .ZN(n4277) );
  NAND2_X1 U35450 ( .A1(n4277), .A2(n2600), .ZN(n2866) );
  NAND2_X1 U35460 ( .A1(n3895), .A2(REG0_REG_22__SCAN_IN), .ZN(n2865) );
  NAND2_X1 U35470 ( .A1(n2598), .A2(REG1_REG_22__SCAN_IN), .ZN(n2864) );
  NAND2_X1 U35480 ( .A1(n2840), .A2(REG2_REG_22__SCAN_IN), .ZN(n2863) );
  OAI22_X1 U35490 ( .A1(n4288), .A2(n2946), .B1(n2945), .B2(n4276), .ZN(n2867)
         );
  XNOR2_X1 U35500 ( .A(n2867), .B(n2233), .ZN(n2871) );
  OR2_X1 U35510 ( .A1(n4288), .A2(n2947), .ZN(n2869) );
  NAND2_X1 U35520 ( .A1(n2913), .A2(n3046), .ZN(n2868) );
  NAND2_X1 U35530 ( .A1(n2869), .A2(n2868), .ZN(n2870) );
  XNOR2_X1 U35540 ( .A(n2871), .B(n2870), .ZN(n3821) );
  NOR2_X1 U35550 ( .A1(n2871), .A2(n2870), .ZN(n3663) );
  INV_X1 U35560 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4433) );
  INV_X1 U35570 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3822) );
  INV_X1 U35580 ( .A(REG3_REG_23__SCAN_IN), .ZN(n5072) );
  OAI21_X1 U35590 ( .B1(n2873), .B2(n3822), .A(n5072), .ZN(n2874) );
  NAND2_X1 U35600 ( .A1(REG3_REG_23__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2872) );
  AND2_X1 U35610 ( .A1(n2874), .A2(n2885), .ZN(n4263) );
  NAND2_X1 U35620 ( .A1(n4263), .A2(n2600), .ZN(n2878) );
  NAND2_X1 U35630 ( .A1(n2840), .A2(REG2_REG_23__SCAN_IN), .ZN(n2876) );
  NAND2_X1 U35640 ( .A1(n3895), .A2(REG0_REG_23__SCAN_IN), .ZN(n2875) );
  AND2_X1 U35650 ( .A1(n2876), .A2(n2875), .ZN(n2877) );
  OAI211_X1 U35660 ( .C1(n2564), .C2(n4433), .A(n2878), .B(n2877), .ZN(n4054)
         );
  NAND2_X1 U35670 ( .A1(n4054), .A2(n2984), .ZN(n2880) );
  NAND2_X1 U35680 ( .A1(n2914), .A2(n4260), .ZN(n2879) );
  NAND2_X1 U35690 ( .A1(n2880), .A2(n2879), .ZN(n2881) );
  XNOR2_X1 U35700 ( .A(n2881), .B(n2917), .ZN(n2884) );
  NOR2_X1 U35710 ( .A1(n2946), .A2(n4254), .ZN(n2882) );
  AOI21_X1 U35720 ( .B1(n4054), .B2(n2920), .A(n2882), .ZN(n2883) );
  XNOR2_X1 U35730 ( .A(n2884), .B(n2883), .ZN(n3662) );
  AND2_X1 U35740 ( .A1(n2885), .A2(n4975), .ZN(n2886) );
  OR2_X1 U35750 ( .A1(n2886), .A2(n2907), .ZN(n3771) );
  AOI22_X1 U35760 ( .A1(n2840), .A2(REG2_REG_24__SCAN_IN), .B1(n3895), .B2(
        REG0_REG_24__SCAN_IN), .ZN(n2889) );
  NAND2_X1 U35770 ( .A1(n2598), .A2(REG1_REG_24__SCAN_IN), .ZN(n2888) );
  NAND2_X1 U35780 ( .A1(n4212), .A2(n2920), .ZN(n2891) );
  NAND2_X1 U35790 ( .A1(n2984), .A2(n4237), .ZN(n2890) );
  INV_X1 U35800 ( .A(n4212), .ZN(n4255) );
  OAI22_X1 U35810 ( .A1(n4255), .A2(n2946), .B1(n2945), .B2(n4424), .ZN(n2893)
         );
  XOR2_X1 U3582 ( .A(n2234), .B(n2893), .Z(n3768) );
  INV_X1 U3583 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4879) );
  XNOR2_X1 U3584 ( .A(n2907), .B(n4879), .ZN(n4221) );
  NAND2_X1 U3585 ( .A1(n4221), .A2(n2600), .ZN(n2898) );
  INV_X1 U3586 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4422) );
  NAND2_X1 U3587 ( .A1(n2840), .A2(REG2_REG_25__SCAN_IN), .ZN(n2895) );
  NAND2_X1 U3588 ( .A1(n3895), .A2(REG0_REG_25__SCAN_IN), .ZN(n2894) );
  OAI211_X1 U3589 ( .C1(n4422), .C2(n2564), .A(n2895), .B(n2894), .ZN(n2896)
         );
  INV_X1 U3590 ( .A(n2896), .ZN(n2897) );
  NAND2_X1 U3591 ( .A1(n4192), .A2(n2984), .ZN(n2901) );
  NAND2_X1 U3592 ( .A1(n2899), .A2(n4211), .ZN(n2900) );
  NAND2_X1 U3593 ( .A1(n2901), .A2(n2900), .ZN(n2902) );
  XNOR2_X1 U3594 ( .A(n2902), .B(n2917), .ZN(n2905) );
  NOR2_X1 U3595 ( .A1(n2946), .A2(n4219), .ZN(n2903) );
  AOI21_X1 U3596 ( .B1(n4192), .B2(n2920), .A(n2903), .ZN(n2904) );
  NAND2_X1 U3597 ( .A1(n2905), .A2(n2904), .ZN(n3727) );
  NOR2_X1 U3598 ( .A1(n2905), .A2(n2904), .ZN(n3726) );
  AOI21_X2 U3599 ( .B1(n3730), .B2(n3727), .A(n3726), .ZN(n3870) );
  AND2_X1 U3600 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2906) );
  AOI21_X1 U3601 ( .B1(n2907), .B2(REG3_REG_25__SCAN_IN), .A(
        REG3_REG_26__SCAN_IN), .ZN(n2908) );
  INV_X1 U3602 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4418) );
  NAND2_X1 U3603 ( .A1(n2840), .A2(REG2_REG_26__SCAN_IN), .ZN(n2910) );
  NAND2_X1 U3604 ( .A1(n3895), .A2(REG0_REG_26__SCAN_IN), .ZN(n2909) );
  OAI211_X1 U3605 ( .C1(n4418), .C2(n2564), .A(n2910), .B(n2909), .ZN(n2911)
         );
  INV_X1 U3606 ( .A(n2911), .ZN(n2912) );
  NAND2_X1 U3607 ( .A1(n4409), .A2(n2913), .ZN(n2916) );
  NAND2_X1 U3608 ( .A1(n2914), .A2(n3872), .ZN(n2915) );
  NAND2_X1 U3609 ( .A1(n2916), .A2(n2915), .ZN(n2918) );
  XNOR2_X1 U3610 ( .A(n2918), .B(n2917), .ZN(n2924) );
  INV_X1 U3611 ( .A(n2924), .ZN(n2922) );
  NOR2_X1 U3612 ( .A1(n2946), .A2(n4199), .ZN(n2919) );
  AOI21_X1 U3613 ( .B1(n4409), .B2(n2920), .A(n2919), .ZN(n2923) );
  INV_X1 U3614 ( .A(n2923), .ZN(n2921) );
  NAND2_X1 U3615 ( .A1(n2922), .A2(n2921), .ZN(n3867) );
  AND2_X1 U3616 ( .A1(n2924), .A2(n2923), .ZN(n3868) );
  NAND2_X1 U3617 ( .A1(n2925), .A2(REG3_REG_27__SCAN_IN), .ZN(n2937) );
  OR2_X1 U3618 ( .A1(n2925), .A2(REG3_REG_27__SCAN_IN), .ZN(n2926) );
  NAND2_X1 U3619 ( .A1(n4173), .A2(n2600), .ZN(n2932) );
  INV_X1 U3620 ( .A(REG1_REG_27__SCAN_IN), .ZN(n2929) );
  NAND2_X1 U3621 ( .A1(n2840), .A2(REG2_REG_27__SCAN_IN), .ZN(n2928) );
  NAND2_X1 U3622 ( .A1(n3895), .A2(REG0_REG_27__SCAN_IN), .ZN(n2927) );
  OAI211_X1 U3623 ( .C1(n2929), .C2(n2564), .A(n2928), .B(n2927), .ZN(n2930)
         );
  INV_X1 U3624 ( .A(n2930), .ZN(n2931) );
  OAI22_X1 U3625 ( .A1(n4185), .A2(n2947), .B1(n4170), .B2(n2933), .ZN(n2935)
         );
  OAI22_X1 U3626 ( .A1(n4185), .A2(n2946), .B1(n4170), .B2(n2945), .ZN(n2934)
         );
  XNOR2_X1 U3627 ( .A(n2934), .B(n2234), .ZN(n2936) );
  NAND2_X1 U3628 ( .A1(n2937), .A2(n4846), .ZN(n2938) );
  NAND2_X1 U3629 ( .A1(n3626), .A2(n2938), .ZN(n2988) );
  INV_X1 U3630 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2941) );
  NAND2_X1 U3631 ( .A1(n2840), .A2(REG2_REG_28__SCAN_IN), .ZN(n2940) );
  NAND2_X1 U3632 ( .A1(n3895), .A2(REG0_REG_28__SCAN_IN), .ZN(n2939) );
  OAI211_X1 U3633 ( .C1(n2941), .C2(n2564), .A(n2940), .B(n2939), .ZN(n2942)
         );
  INV_X1 U3634 ( .A(n2942), .ZN(n2943) );
  INV_X1 U3635 ( .A(n4179), .ZN(n3624) );
  OAI22_X1 U3636 ( .A1(n3624), .A2(n2946), .B1(n2945), .B2(n4157), .ZN(n2951)
         );
  OAI22_X1 U3637 ( .A1(n3624), .A2(n2947), .B1(n2946), .B2(n4157), .ZN(n2949)
         );
  XNOR2_X1 U3638 ( .A(n2949), .B(n2233), .ZN(n2950) );
  XOR2_X1 U3639 ( .A(n2951), .B(n2950), .Z(n2952) );
  NAND2_X1 U3640 ( .A1(n3116), .A2(B_REG_SCAN_IN), .ZN(n2954) );
  MUX2_X1 U3641 ( .A(n2954), .B(B_REG_SCAN_IN), .S(n2953), .Z(n2955) );
  INV_X1 U3642 ( .A(n2953), .ZN(n2956) );
  NAND2_X1 U3643 ( .A1(n2956), .A2(n2969), .ZN(n3139) );
  NOR4_X1 U3644 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2961) );
  NOR4_X1 U3645 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n2960) );
  NOR4_X1 U3646 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2959) );
  NOR4_X1 U3647 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2958) );
  NAND4_X1 U3648 ( .A1(n2961), .A2(n2960), .A3(n2959), .A4(n2958), .ZN(n2967)
         );
  NOR2_X1 U3649 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_27__SCAN_IN), .ZN(n2965)
         );
  NOR4_X1 U3650 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2964) );
  NOR4_X1 U3651 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2963) );
  NOR4_X1 U3652 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2962) );
  NAND4_X1 U3653 ( .A1(n2965), .A2(n2964), .A3(n2963), .A4(n2962), .ZN(n2966)
         );
  NOR2_X1 U3654 ( .A1(n2967), .A2(n2966), .ZN(n2968) );
  NAND2_X1 U3655 ( .A1(n2969), .A2(n3116), .ZN(n3137) );
  NAND2_X1 U3656 ( .A1(n2506), .A2(n4144), .ZN(n2978) );
  NAND2_X1 U3657 ( .A1(n3311), .A2(n2978), .ZN(n2973) );
  AND2_X1 U3658 ( .A1(n4048), .A2(n4539), .ZN(n3131) );
  INV_X1 U3659 ( .A(n3131), .ZN(n2972) );
  NAND2_X1 U3660 ( .A1(n2973), .A2(n2972), .ZN(n2976) );
  NOR2_X1 U3661 ( .A1(n3275), .A2(n2976), .ZN(n2974) );
  INV_X1 U3662 ( .A(n3007), .ZN(n2986) );
  OR2_X2 U3663 ( .A1(n2975), .A2(n2506), .ZN(n4459) );
  NAND2_X1 U3664 ( .A1(n2976), .A2(n4459), .ZN(n2977) );
  NAND2_X1 U3665 ( .A1(n2986), .A2(n2977), .ZN(n2979) );
  NAND2_X1 U3666 ( .A1(n3131), .A2(n2978), .ZN(n3277) );
  NAND2_X1 U3667 ( .A1(n2979), .A2(n3277), .ZN(n3231) );
  NAND2_X1 U3668 ( .A1(n2536), .A2(n3132), .ZN(n2980) );
  OAI21_X1 U3669 ( .B1(n3231), .B2(n2980), .A(STATE_REG_SCAN_IN), .ZN(n2987)
         );
  INV_X1 U3670 ( .A(n2981), .ZN(n2982) );
  AND2_X1 U3671 ( .A1(n4660), .A2(n2982), .ZN(n2983) );
  NAND2_X1 U3672 ( .A1(n2984), .A2(n2983), .ZN(n4047) );
  INV_X1 U3673 ( .A(n4047), .ZN(n2985) );
  NAND2_X1 U3674 ( .A1(n2986), .A2(n2985), .ZN(n3232) );
  INV_X1 U3675 ( .A(n2988), .ZN(n4158) );
  NAND2_X1 U3676 ( .A1(n3890), .A2(n4158), .ZN(n3012) );
  INV_X1 U3677 ( .A(n4185), .ZN(n4400) );
  NAND2_X1 U3678 ( .A1(n2989), .A2(IR_REG_31__SCAN_IN), .ZN(n2990) );
  MUX2_X1 U3679 ( .A(n2990), .B(IR_REG_31__SCAN_IN), .S(n2436), .Z(n2992) );
  NAND2_X1 U3680 ( .A1(n2992), .A2(n2468), .ZN(n3189) );
  NOR2_X1 U3681 ( .A1(n4047), .A2(n3189), .ZN(n2993) );
  AND2_X2 U3682 ( .A1(n3007), .A2(n2993), .ZN(n3886) );
  NOR2_X1 U3683 ( .A1(n3275), .A2(n4459), .ZN(n2994) );
  NAND2_X1 U3684 ( .A1(n3007), .A2(n2994), .ZN(n2998) );
  AND2_X1 U3685 ( .A1(n2506), .A2(n4540), .ZN(n3314) );
  AND2_X1 U3686 ( .A1(n3314), .A2(n2995), .ZN(n4699) );
  NAND2_X1 U3687 ( .A1(n4699), .A2(n2996), .ZN(n3101) );
  INV_X2 U3688 ( .A(n3825), .ZN(n3887) );
  AOI22_X1 U3689 ( .A1(n4400), .A2(n3886), .B1(n2324), .B2(n3887), .ZN(n3010)
         );
  INV_X1 U3690 ( .A(n3626), .ZN(n2999) );
  NAND2_X1 U3691 ( .A1(n2999), .A2(n2600), .ZN(n3005) );
  INV_X1 U3692 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3002) );
  NAND2_X1 U3693 ( .A1(n2840), .A2(REG2_REG_29__SCAN_IN), .ZN(n3001) );
  NAND2_X1 U3694 ( .A1(n3895), .A2(REG0_REG_29__SCAN_IN), .ZN(n3000) );
  OAI211_X1 U3695 ( .C1(n2564), .C2(n3002), .A(n3001), .B(n3000), .ZN(n3003)
         );
  INV_X1 U3696 ( .A(n3003), .ZN(n3004) );
  NAND2_X1 U3697 ( .A1(n3005), .A2(n3004), .ZN(n4163) );
  INV_X1 U3698 ( .A(n3189), .ZN(n3148) );
  NOR2_X1 U3699 ( .A1(n4047), .A2(n3148), .ZN(n3006) );
  AND2_X2 U3700 ( .A1(n3007), .A2(n3006), .ZN(n3885) );
  NOR2_X1 U3701 ( .A1(n4846), .A2(STATE_REG_SCAN_IN), .ZN(n3008) );
  AOI21_X1 U3702 ( .B1(n4163), .B2(n3885), .A(n3008), .ZN(n3009) );
  NAND2_X1 U3703 ( .A1(n3014), .A2(n3013), .ZN(U3217) );
  INV_X1 U3704 ( .A(n2557), .ZN(n3015) );
  AND2_X1 U3705 ( .A1(n4072), .A2(n3312), .ZN(n3281) );
  NAND2_X1 U3706 ( .A1(n3056), .A2(n3281), .ZN(n3283) );
  NAND2_X1 U3707 ( .A1(n4070), .A2(n3241), .ZN(n3016) );
  NAND2_X1 U3708 ( .A1(n3283), .A2(n3016), .ZN(n3321) );
  INV_X1 U3709 ( .A(n3321), .ZN(n3018) );
  NAND2_X1 U3710 ( .A1(n3017), .A2(n3106), .ZN(n3936) );
  NAND2_X1 U3711 ( .A1(n2574), .A2(n3330), .ZN(n3939) );
  NAND2_X1 U3712 ( .A1(n3018), .A2(n3057), .ZN(n3319) );
  NAND2_X1 U3713 ( .A1(n3017), .A2(n3330), .ZN(n3019) );
  NAND2_X1 U3714 ( .A1(n3319), .A2(n3019), .ZN(n3265) );
  NOR2_X1 U3715 ( .A1(n2592), .A2(n3262), .ZN(n3020) );
  INV_X1 U3716 ( .A(n2592), .ZN(n3302) );
  OAI22_X1 U3717 ( .A1(n3265), .A2(n3020), .B1(n3302), .B2(n3395), .ZN(n3299)
         );
  INV_X1 U3718 ( .A(n4069), .ZN(n3385) );
  NAND2_X1 U3719 ( .A1(n4069), .A2(n3297), .ZN(n3945) );
  NAND2_X1 U3720 ( .A1(n3942), .A2(n3945), .ZN(n3910) );
  NAND2_X1 U3721 ( .A1(n3299), .A2(n3910), .ZN(n3022) );
  NAND2_X1 U3722 ( .A1(n4069), .A2(n3781), .ZN(n3021) );
  NAND2_X1 U3723 ( .A1(n3022), .A2(n3021), .ZN(n3337) );
  AND2_X1 U3724 ( .A1(n4068), .A2(n3749), .ZN(n3024) );
  INV_X1 U3725 ( .A(n4068), .ZN(n3404) );
  NAND2_X1 U3726 ( .A1(n3404), .A2(n3339), .ZN(n3023) );
  NOR2_X1 U3727 ( .A1(n4067), .A2(n3861), .ZN(n3025) );
  INV_X1 U3728 ( .A(n4066), .ZN(n3475) );
  NAND2_X1 U3729 ( .A1(n3475), .A2(n3638), .ZN(n3062) );
  NAND2_X1 U3730 ( .A1(n4066), .A2(n3360), .ZN(n3951) );
  NAND2_X1 U3731 ( .A1(n3062), .A2(n3951), .ZN(n3920) );
  AND2_X1 U3732 ( .A1(n4065), .A2(n3696), .ZN(n3026) );
  OAI22_X1 U3733 ( .A1(n3472), .A2(n3026), .B1(n3696), .B2(n4065), .ZN(n3415)
         );
  NAND2_X1 U3734 ( .A1(n4064), .A2(n3790), .ZN(n3027) );
  AND2_X1 U3735 ( .A1(n4063), .A2(n3674), .ZN(n3029) );
  INV_X1 U3736 ( .A(n4063), .ZN(n3413) );
  NAND2_X1 U3737 ( .A1(n3413), .A2(n3534), .ZN(n3028) );
  INV_X1 U3738 ( .A(n4062), .ZN(n3547) );
  NAND2_X1 U3739 ( .A1(n3547), .A2(n3837), .ZN(n3485) );
  NAND2_X1 U3740 ( .A1(n4062), .A2(n3508), .ZN(n3487) );
  NAND2_X1 U3741 ( .A1(n3485), .A2(n3487), .ZN(n3921) );
  NAND2_X1 U3742 ( .A1(n3501), .A2(n3921), .ZN(n3031) );
  NAND2_X1 U3743 ( .A1(n3547), .A2(n3508), .ZN(n3030) );
  NAND2_X1 U3744 ( .A1(n3031), .A2(n3030), .ZN(n3489) );
  NOR2_X1 U3745 ( .A1(n4061), .A2(n3720), .ZN(n3032) );
  INV_X1 U3746 ( .A(n4061), .ZN(n3502) );
  INV_X1 U3747 ( .A(n3720), .ZN(n3546) );
  AND2_X1 U3748 ( .A1(n4060), .A2(n3813), .ZN(n3034) );
  NAND2_X1 U3749 ( .A1(n3577), .A2(n3518), .ZN(n3033) );
  NAND2_X1 U3750 ( .A1(n3595), .A2(n3656), .ZN(n3977) );
  NAND2_X1 U3751 ( .A1(n4059), .A2(n3581), .ZN(n3957) );
  NAND2_X1 U3752 ( .A1(n3977), .A2(n3957), .ZN(n3906) );
  NAND2_X1 U3753 ( .A1(n3595), .A2(n3581), .ZN(n3035) );
  NAND2_X1 U3754 ( .A1(n4058), .A2(n3888), .ZN(n3036) );
  NAND2_X1 U3755 ( .A1(n3037), .A2(n3036), .ZN(n3606) );
  NAND2_X1 U3756 ( .A1(n4461), .A2(n3739), .ZN(n4013) );
  NAND2_X1 U3757 ( .A1(n4057), .A2(n3617), .ZN(n3979) );
  NAND2_X1 U3758 ( .A1(n4013), .A2(n3979), .ZN(n3613) );
  NAND2_X1 U3759 ( .A1(n3606), .A2(n3613), .ZN(n3605) );
  NAND2_X1 U3760 ( .A1(n3605), .A2(n2446), .ZN(n4364) );
  INV_X1 U3761 ( .A(n4056), .ZN(n4352) );
  NAND2_X1 U3762 ( .A1(n4352), .A2(n4458), .ZN(n3039) );
  AOI21_X1 U3763 ( .B1(n4364), .B2(n3039), .A(n3038), .ZN(n4345) );
  INV_X1 U3764 ( .A(n4370), .ZN(n3040) );
  NAND2_X1 U3765 ( .A1(n3040), .A2(n4349), .ZN(n4326) );
  NAND2_X1 U3766 ( .A1(n4370), .A2(n4357), .ZN(n4327) );
  NAND2_X1 U3767 ( .A1(n4326), .A2(n4327), .ZN(n4348) );
  NAND2_X1 U3768 ( .A1(n4055), .A2(n4306), .ZN(n3913) );
  NOR2_X1 U3769 ( .A1(n4055), .A2(n4306), .ZN(n3914) );
  AOI21_X2 U3770 ( .B1(n4301), .B2(n3913), .A(n3914), .ZN(n4283) );
  INV_X1 U3771 ( .A(n4288), .ZN(n4257) );
  NAND2_X1 U3772 ( .A1(n4257), .A2(n4276), .ZN(n3084) );
  NAND2_X1 U3773 ( .A1(n4288), .A2(n3046), .ZN(n4251) );
  NAND2_X1 U3774 ( .A1(n3084), .A2(n4251), .ZN(n4271) );
  NAND2_X1 U3775 ( .A1(n4425), .A2(n4254), .ZN(n3048) );
  NAND2_X1 U3776 ( .A1(n4212), .A2(n4237), .ZN(n3050) );
  NAND2_X1 U3777 ( .A1(n4206), .A2(n3051), .ZN(n3052) );
  INV_X1 U3778 ( .A(n4192), .ZN(n4231) );
  NAND2_X1 U3779 ( .A1(n3052), .A2(n2452), .ZN(n4193) );
  NOR2_X1 U3780 ( .A1(n4409), .A2(n3872), .ZN(n3053) );
  NOR2_X1 U3781 ( .A1(n4179), .A2(n4157), .ZN(n4029) );
  NAND2_X1 U3782 ( .A1(n2552), .A2(DATAI_29_), .ZN(n3107) );
  XNOR2_X1 U3783 ( .A(n4163), .B(n3107), .ZN(n3899) );
  XNOR2_X1 U3784 ( .A(n3054), .B(n3899), .ZN(n3622) );
  XNOR2_X1 U3785 ( .A(n2507), .B(n4048), .ZN(n3055) );
  NAND2_X1 U3786 ( .A1(n3055), .A2(n4144), .ZN(n4312) );
  INV_X1 U3787 ( .A(n4699), .ZN(n4674) );
  NOR2_X1 U3788 ( .A1(n4459), .A2(n3107), .ZN(n3099) );
  INV_X1 U3789 ( .A(n4072), .ZN(n3239) );
  NAND2_X1 U3790 ( .A1(n3239), .A2(n3312), .ZN(n3931) );
  NAND2_X1 U3791 ( .A1(n3318), .A2(n3320), .ZN(n3058) );
  NAND2_X1 U3792 ( .A1(n3058), .A2(n3936), .ZN(n3267) );
  NAND2_X1 U3793 ( .A1(n3302), .A2(n3262), .ZN(n3941) );
  NAND2_X1 U3794 ( .A1(n2592), .A2(n3395), .ZN(n3938) );
  AND2_X1 U3795 ( .A1(n3941), .A2(n3938), .ZN(n3266) );
  NAND2_X1 U3796 ( .A1(n3267), .A2(n3266), .ZN(n3059) );
  INV_X1 U3797 ( .A(n3942), .ZN(n3060) );
  AND2_X1 U3798 ( .A1(n4068), .A2(n3339), .ZN(n3338) );
  NAND2_X1 U3799 ( .A1(n3404), .A2(n3749), .ZN(n3961) );
  NAND2_X1 U3800 ( .A1(n4067), .A2(n3370), .ZN(n3959) );
  NAND2_X1 U3801 ( .A1(n3367), .A2(n3959), .ZN(n3061) );
  INV_X1 U3802 ( .A(n4067), .ZN(n3341) );
  NAND2_X1 U3803 ( .A1(n3341), .A2(n3861), .ZN(n3947) );
  NAND2_X1 U3804 ( .A1(n3061), .A2(n3947), .ZN(n3352) );
  INV_X1 U3805 ( .A(n3062), .ZN(n3063) );
  OR2_X1 U3806 ( .A1(n3352), .A2(n3063), .ZN(n3064) );
  NAND2_X1 U3807 ( .A1(n3064), .A2(n3951), .ZN(n3473) );
  INV_X1 U3808 ( .A(n4065), .ZN(n3460) );
  NAND2_X1 U3809 ( .A1(n3460), .A2(n3696), .ZN(n3953) );
  INV_X1 U3810 ( .A(n3696), .ZN(n3474) );
  NAND2_X1 U3811 ( .A1(n4065), .A2(n3474), .ZN(n3950) );
  AND2_X1 U3812 ( .A1(n4064), .A2(n3459), .ZN(n3969) );
  INV_X1 U3813 ( .A(n4064), .ZN(n3535) );
  NAND2_X1 U3814 ( .A1(n3535), .A2(n3790), .ZN(n3952) );
  NAND2_X1 U3815 ( .A1(n4063), .A2(n3534), .ZN(n3972) );
  NAND2_X1 U3816 ( .A1(n3533), .A2(n3972), .ZN(n3065) );
  NAND2_X1 U3817 ( .A1(n3413), .A2(n3674), .ZN(n3970) );
  NAND2_X1 U3818 ( .A1(n3065), .A2(n3970), .ZN(n3500) );
  NAND2_X1 U3819 ( .A1(n4061), .A2(n3546), .ZN(n3513) );
  NAND2_X1 U3820 ( .A1(n4060), .A2(n3518), .ZN(n3066) );
  NAND2_X1 U3821 ( .A1(n3513), .A2(n3066), .ZN(n3068) );
  INV_X1 U3822 ( .A(n3487), .ZN(n3067) );
  NOR2_X1 U3823 ( .A1(n3068), .A2(n3067), .ZN(n3973) );
  NAND2_X1 U3824 ( .A1(n3500), .A2(n3973), .ZN(n3072) );
  NAND2_X1 U3825 ( .A1(n3502), .A2(n3720), .ZN(n3515) );
  NAND2_X1 U3826 ( .A1(n3485), .A2(n3515), .ZN(n3071) );
  INV_X1 U3827 ( .A(n3068), .ZN(n3070) );
  NOR2_X1 U3828 ( .A1(n4060), .A2(n3518), .ZN(n3069) );
  AOI21_X1 U3829 ( .B1(n3071), .B2(n3070), .A(n3069), .ZN(n3975) );
  NAND2_X1 U3830 ( .A1(n3072), .A2(n3975), .ZN(n4011) );
  INV_X1 U3831 ( .A(n3906), .ZN(n3573) );
  NAND2_X1 U3832 ( .A1(n3073), .A2(n3888), .ZN(n3976) );
  NAND2_X1 U3833 ( .A1(n4058), .A2(n3594), .ZN(n3958) );
  NAND2_X1 U3834 ( .A1(n3976), .A2(n3958), .ZN(n3905) );
  INV_X1 U3835 ( .A(n3977), .ZN(n3074) );
  NOR2_X1 U3836 ( .A1(n3905), .A2(n3074), .ZN(n3075) );
  INV_X1 U3837 ( .A(n3613), .ZN(n3904) );
  NAND2_X1 U3838 ( .A1(n3076), .A2(n3979), .ZN(n4366) );
  NAND2_X1 U3839 ( .A1(n4352), .A2(n4383), .ZN(n4324) );
  NAND2_X1 U3840 ( .A1(n4326), .A2(n4324), .ZN(n3079) );
  NAND2_X1 U3841 ( .A1(n4350), .A2(n4336), .ZN(n3077) );
  AND2_X1 U3842 ( .A1(n4327), .A2(n3077), .ZN(n4246) );
  NOR2_X1 U3843 ( .A1(n4350), .A2(n4336), .ZN(n3078) );
  AOI21_X1 U3844 ( .B1(n3079), .B2(n4246), .A(n3078), .ZN(n4302) );
  INV_X1 U3845 ( .A(n4055), .ZN(n4441) );
  NAND2_X1 U3846 ( .A1(n4441), .A2(n4306), .ZN(n3080) );
  NAND2_X1 U3847 ( .A1(n4366), .A2(n4249), .ZN(n3081) );
  NAND2_X1 U3848 ( .A1(n4056), .A2(n4458), .ZN(n4244) );
  NAND2_X1 U3849 ( .A1(n4246), .A2(n4244), .ZN(n3982) );
  AND2_X1 U3850 ( .A1(n4055), .A2(n4314), .ZN(n4248) );
  AOI21_X1 U3851 ( .B1(n4249), .B2(n3982), .A(n4248), .ZN(n4015) );
  NAND2_X1 U3852 ( .A1(n3081), .A2(n4015), .ZN(n3083) );
  NAND2_X1 U3853 ( .A1(n4308), .A2(n4296), .ZN(n4250) );
  NAND2_X1 U3854 ( .A1(n4251), .A2(n4250), .ZN(n4020) );
  INV_X1 U3855 ( .A(n4020), .ZN(n3082) );
  NAND2_X1 U3856 ( .A1(n3083), .A2(n3082), .ZN(n3088) );
  NAND2_X1 U3857 ( .A1(n4054), .A2(n4254), .ZN(n3085) );
  NAND2_X1 U3858 ( .A1(n3085), .A2(n3084), .ZN(n3989) );
  INV_X1 U3859 ( .A(n3989), .ZN(n3087) );
  AND2_X1 U3860 ( .A1(n4273), .A2(n4440), .ZN(n3986) );
  NAND2_X1 U3861 ( .A1(n4251), .A2(n3986), .ZN(n3086) );
  AND2_X1 U3862 ( .A1(n3087), .A2(n3086), .ZN(n4019) );
  OR2_X1 U3863 ( .A1(n4212), .A2(n4424), .ZN(n3912) );
  NAND2_X1 U3864 ( .A1(n4425), .A2(n4260), .ZN(n4227) );
  NAND2_X1 U3865 ( .A1(n4192), .A2(n4219), .ZN(n3930) );
  NOR2_X1 U3866 ( .A1(n4409), .A2(n4199), .ZN(n3900) );
  NOR2_X1 U3867 ( .A1(n4192), .A2(n4219), .ZN(n4186) );
  NOR2_X1 U3868 ( .A1(n3900), .A2(n4186), .ZN(n4022) );
  AND2_X1 U3869 ( .A1(n4409), .A2(n4199), .ZN(n3993) );
  NOR2_X1 U3870 ( .A1(n4185), .A2(n4407), .ZN(n3995) );
  INV_X1 U3871 ( .A(n4028), .ZN(n3089) );
  OAI21_X1 U3872 ( .B1(n4178), .B2(n4177), .A(n3089), .ZN(n4162) );
  INV_X1 U3873 ( .A(n3090), .ZN(n3992) );
  AOI21_X1 U3874 ( .B1(n4162), .B2(n3992), .A(n4029), .ZN(n3091) );
  XOR2_X1 U3875 ( .A(n3899), .B(n3091), .Z(n3098) );
  INV_X1 U3876 ( .A(n2506), .ZN(n4005) );
  NAND2_X1 U3877 ( .A1(n4005), .A2(n4539), .ZN(n4038) );
  NAND2_X1 U3878 ( .A1(n4048), .A2(n4540), .ZN(n3092) );
  NAND2_X1 U3879 ( .A1(n2840), .A2(REG2_REG_30__SCAN_IN), .ZN(n3094) );
  NAND2_X1 U3880 ( .A1(n3895), .A2(REG0_REG_30__SCAN_IN), .ZN(n3093) );
  OAI211_X1 U3881 ( .C1(n2564), .C2(n4398), .A(n3094), .B(n3093), .ZN(n4053)
         );
  INV_X1 U3882 ( .A(n4053), .ZN(n3097) );
  XNOR2_X1 U3883 ( .A(n3095), .B(IR_REG_27__SCAN_IN), .ZN(n3191) );
  NAND2_X1 U3884 ( .A1(n3191), .A2(B_REG_SCAN_IN), .ZN(n3096) );
  NAND2_X1 U3885 ( .A1(n4369), .A2(n3096), .ZN(n4149) );
  OAI22_X1 U3886 ( .A1(n3098), .A2(n4334), .B1(n3097), .B2(n4149), .ZN(n3629)
         );
  NAND2_X1 U3887 ( .A1(n3100), .A2(n3137), .ZN(n3105) );
  NAND2_X1 U3888 ( .A1(n3101), .A2(n3277), .ZN(n3102) );
  NOR2_X1 U3889 ( .A1(n3102), .A2(n3275), .ZN(n3104) );
  NAND3_X1 U3890 ( .A1(n3105), .A2(n3104), .A3(n3103), .ZN(n3110) );
  NAND2_X1 U3891 ( .A1(n2247), .A2(n3360), .ZN(n3469) );
  INV_X1 U3892 ( .A(n3107), .ZN(n4000) );
  NAND2_X1 U3893 ( .A1(n3108), .A2(n2454), .ZN(U3547) );
  INV_X1 U3894 ( .A(n3112), .ZN(n3113) );
  NAND2_X1 U3895 ( .A1(n3113), .A2(n2453), .ZN(U3515) );
  INV_X1 U3896 ( .A(n4660), .ZN(n3114) );
  INV_X2 U3897 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U3898 ( .A1(U3149), .A2(DATAI_25_), .ZN(n3115) );
  OAI21_X1 U3899 ( .B1(n3116), .B2(U3149), .A(n3115), .ZN(U3327) );
  INV_X1 U3900 ( .A(DATAI_18_), .ZN(n4977) );
  NAND2_X1 U3901 ( .A1(n4138), .A2(STATE_REG_SCAN_IN), .ZN(n3117) );
  OAI21_X1 U3902 ( .B1(STATE_REG_SCAN_IN), .B2(n4977), .A(n3117), .ZN(U3334)
         );
  INV_X1 U3903 ( .A(DATAI_26_), .ZN(n3120) );
  NAND2_X1 U3904 ( .A1(n3118), .A2(STATE_REG_SCAN_IN), .ZN(n3119) );
  OAI21_X1 U3905 ( .B1(STATE_REG_SCAN_IN), .B2(n3120), .A(n3119), .ZN(U3326)
         );
  INV_X1 U3906 ( .A(DATAI_27_), .ZN(n4843) );
  NAND2_X1 U3907 ( .A1(n3191), .A2(STATE_REG_SCAN_IN), .ZN(n3121) );
  OAI21_X1 U3908 ( .B1(STATE_REG_SCAN_IN), .B2(n4843), .A(n3121), .ZN(U3325)
         );
  INV_X1 U3909 ( .A(DATAI_20_), .ZN(n3123) );
  NAND2_X1 U3910 ( .A1(n4005), .A2(STATE_REG_SCAN_IN), .ZN(n3122) );
  OAI21_X1 U3911 ( .B1(STATE_REG_SCAN_IN), .B2(n3123), .A(n3122), .ZN(U3332)
         );
  INV_X1 U3912 ( .A(DATAI_22_), .ZN(n4866) );
  NAND2_X1 U3913 ( .A1(n4048), .A2(STATE_REG_SCAN_IN), .ZN(n3124) );
  OAI21_X1 U3914 ( .B1(STATE_REG_SCAN_IN), .B2(n4866), .A(n3124), .ZN(U3330)
         );
  INV_X1 U3915 ( .A(DATAI_24_), .ZN(n3126) );
  NAND2_X1 U3916 ( .A1(n2953), .A2(STATE_REG_SCAN_IN), .ZN(n3125) );
  OAI21_X1 U3917 ( .B1(STATE_REG_SCAN_IN), .B2(n3126), .A(n3125), .ZN(U3328)
         );
  INV_X1 U3918 ( .A(DATAI_30_), .ZN(n3129) );
  NAND2_X1 U3919 ( .A1(n3127), .A2(STATE_REG_SCAN_IN), .ZN(n3128) );
  OAI21_X1 U3920 ( .B1(STATE_REG_SCAN_IN), .B2(n3129), .A(n3128), .ZN(U3322)
         );
  INV_X1 U3921 ( .A(DATAI_28_), .ZN(n4974) );
  NAND2_X1 U3922 ( .A1(n3148), .A2(STATE_REG_SCAN_IN), .ZN(n3130) );
  OAI21_X1 U3923 ( .B1(STATE_REG_SCAN_IN), .B2(n4974), .A(n3130), .ZN(U3324)
         );
  OR2_X1 U3924 ( .A1(n3132), .A2(U3149), .ZN(n4051) );
  NAND2_X1 U3925 ( .A1(n3275), .A2(n4051), .ZN(n3147) );
  NAND2_X1 U3926 ( .A1(n3132), .A2(n3131), .ZN(n3134) );
  INV_X1 U3927 ( .A(n3146), .ZN(n3135) );
  NOR2_X1 U3928 ( .A1(n4628), .A2(U4043), .ZN(U3148) );
  INV_X1 U3929 ( .A(D_REG_1__SCAN_IN), .ZN(n5070) );
  INV_X1 U3930 ( .A(n3137), .ZN(n3138) );
  AOI22_X1 U3931 ( .A1(n4659), .A2(n5070), .B1(n3138), .B2(n4660), .ZN(U3459)
         );
  INV_X1 U3932 ( .A(D_REG_0__SCAN_IN), .ZN(n5075) );
  INV_X1 U3933 ( .A(n3139), .ZN(n3140) );
  AOI22_X1 U3934 ( .A1(n4659), .A2(n5075), .B1(n3140), .B2(n4660), .ZN(U3458)
         );
  NAND2_X1 U3935 ( .A1(n4549), .A2(REG2_REG_1__SCAN_IN), .ZN(n3199) );
  INV_X1 U3936 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3141) );
  MUX2_X1 U3937 ( .A(REG2_REG_1__SCAN_IN), .B(n3141), .S(n4549), .Z(n4084) );
  INV_X1 U3938 ( .A(n3142), .ZN(n3143) );
  AOI22_X1 U3939 ( .A1(n4096), .A2(REG2_REG_3__SCAN_IN), .B1(n4547), .B2(n3143), .ZN(n3144) );
  XNOR2_X1 U3940 ( .A(n3144), .B(n4546), .ZN(n3209) );
  INV_X1 U3941 ( .A(n3144), .ZN(n3145) );
  INV_X1 U3942 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3380) );
  MUX2_X1 U3943 ( .A(n3380), .B(REG2_REG_5__SCAN_IN), .S(n4545), .Z(n3179) );
  XNOR2_X1 U3944 ( .A(n3168), .B(REG2_REG_6__SCAN_IN), .ZN(n3161) );
  NAND2_X1 U3945 ( .A1(n3148), .A2(n3191), .ZN(n4046) );
  INV_X1 U3946 ( .A(n4046), .ZN(n3149) );
  INV_X1 U3947 ( .A(n4635), .ZN(n4092) );
  AND2_X1 U3948 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3860) );
  AOI21_X1 U3949 ( .B1(n4628), .B2(ADDR_REG_6__SCAN_IN), .A(n3860), .ZN(n3150)
         );
  INV_X1 U3950 ( .A(n3150), .ZN(n3159) );
  MUX2_X1 U3951 ( .A(REG1_REG_2__SCAN_IN), .B(n2563), .S(n4548), .Z(n3197) );
  XNOR2_X1 U3952 ( .A(n4549), .B(n2545), .ZN(n4087) );
  AND2_X1 U3953 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4086)
         );
  NAND2_X1 U3954 ( .A1(n4087), .A2(n4086), .ZN(n4085) );
  NAND2_X1 U3955 ( .A1(n4549), .A2(REG1_REG_1__SCAN_IN), .ZN(n3151) );
  NAND2_X1 U3956 ( .A1(n4085), .A2(n3151), .ZN(n3196) );
  NAND2_X1 U3957 ( .A1(n3197), .A2(n3196), .ZN(n3195) );
  NAND2_X1 U3958 ( .A1(n4548), .A2(REG1_REG_2__SCAN_IN), .ZN(n3152) );
  NAND2_X1 U3959 ( .A1(n3195), .A2(n3152), .ZN(n3154) );
  INV_X1 U3960 ( .A(n4547), .ZN(n3153) );
  XNOR2_X1 U3961 ( .A(n3154), .B(n3153), .ZN(n4094) );
  NAND2_X1 U3962 ( .A1(n4094), .A2(REG1_REG_3__SCAN_IN), .ZN(n4093) );
  NAND2_X1 U3963 ( .A1(n3154), .A2(n4547), .ZN(n3155) );
  NAND2_X1 U3964 ( .A1(n4093), .A2(n3155), .ZN(n3156) );
  INV_X1 U3965 ( .A(n4546), .ZN(n3214) );
  XNOR2_X1 U3966 ( .A(n3156), .B(n3214), .ZN(n3211) );
  XNOR2_X1 U3967 ( .A(n4545), .B(REG1_REG_5__SCAN_IN), .ZN(n3176) );
  NOR2_X1 U3968 ( .A1(n3177), .A2(n3176), .ZN(n3175) );
  AOI21_X1 U3969 ( .B1(REG1_REG_5__SCAN_IN), .B2(n4545), .A(n3175), .ZN(n3162)
         );
  XOR2_X1 U3970 ( .A(n4544), .B(n3162), .Z(n3157) );
  INV_X1 U3971 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3374) );
  INV_X1 U3972 ( .A(n3191), .ZN(n4074) );
  INV_X1 U3973 ( .A(n4629), .ZN(n3174) );
  NOR2_X1 U3974 ( .A1(n3157), .A2(n3374), .ZN(n3163) );
  AOI211_X1 U3975 ( .C1(n3157), .C2(n3374), .A(n3174), .B(n3163), .ZN(n3158)
         );
  AOI211_X1 U3976 ( .C1(n4092), .C2(n4544), .A(n3159), .B(n3158), .ZN(n3160)
         );
  OAI21_X1 U3977 ( .B1(n3161), .B2(n4622), .A(n3160), .ZN(U3246) );
  INV_X1 U3978 ( .A(n4542), .ZN(n3444) );
  INV_X1 U3979 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4708) );
  INV_X1 U3980 ( .A(n4543), .ZN(n3223) );
  XNOR2_X1 U3981 ( .A(n3164), .B(n4542), .ZN(n3428) );
  XNOR2_X1 U3982 ( .A(n3428), .B(REG1_REG_8__SCAN_IN), .ZN(n3165) );
  NAND2_X1 U3983 ( .A1(n3165), .A2(n4629), .ZN(n3173) );
  INV_X1 U3984 ( .A(n3166), .ZN(n3167) );
  INV_X1 U3985 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3362) );
  MUX2_X1 U3986 ( .A(n3362), .B(REG2_REG_7__SCAN_IN), .S(n4543), .Z(n3225) );
  NOR2_X1 U3987 ( .A1(n3226), .A2(n3225), .ZN(n3224) );
  AOI21_X1 U3988 ( .B1(n4543), .B2(REG2_REG_7__SCAN_IN), .A(n3224), .ZN(n3445)
         );
  XNOR2_X1 U3989 ( .A(n3445), .B(n3444), .ZN(n3446) );
  XNOR2_X1 U3990 ( .A(REG2_REG_8__SCAN_IN), .B(n3446), .ZN(n3169) );
  NAND2_X1 U3991 ( .A1(n4587), .A2(n3169), .ZN(n3170) );
  NAND2_X1 U3992 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3694) );
  NAND2_X1 U3993 ( .A1(n3170), .A2(n3694), .ZN(n3171) );
  AOI21_X1 U3994 ( .B1(n4628), .B2(ADDR_REG_8__SCAN_IN), .A(n3171), .ZN(n3172)
         );
  OAI211_X1 U3995 ( .C1(n4635), .C2(n3444), .A(n3173), .B(n3172), .ZN(U3248)
         );
  AOI211_X1 U3996 ( .C1(n3177), .C2(n3176), .A(n3175), .B(n3174), .ZN(n3185)
         );
  AOI211_X1 U3997 ( .C1(n3180), .C2(n3179), .A(n3178), .B(n4622), .ZN(n3184)
         );
  INV_X1 U3998 ( .A(n4545), .ZN(n3182) );
  INV_X1 U3999 ( .A(REG3_REG_5__SCAN_IN), .ZN(n5013) );
  NOR2_X1 U4000 ( .A1(STATE_REG_SCAN_IN), .A2(n5013), .ZN(n3748) );
  AOI21_X1 U4001 ( .B1(n4628), .B2(ADDR_REG_5__SCAN_IN), .A(n3748), .ZN(n3181)
         );
  OAI21_X1 U4002 ( .B1(n4635), .B2(n3182), .A(n3181), .ZN(n3183) );
  OR3_X1 U4003 ( .A1(n3185), .A2(n3184), .A3(n3183), .ZN(U3245) );
  OAI21_X1 U4004 ( .B1(n3188), .B2(n3187), .A(n3186), .ZN(n3235) );
  NOR2_X1 U4005 ( .A1(n3189), .A2(n3191), .ZN(n3193) );
  INV_X1 U4006 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3190) );
  AOI21_X1 U4007 ( .B1(n3191), .B2(n3190), .A(n3189), .ZN(n4073) );
  NAND2_X1 U4008 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4082) );
  OAI22_X1 U4009 ( .A1(n4073), .A2(IR_REG_0__SCAN_IN), .B1(n4082), .B2(n4046), 
        .ZN(n3192) );
  AOI211_X1 U4010 ( .C1(n3235), .C2(n3193), .A(n4071), .B(n3192), .ZN(n3215)
         );
  INV_X1 U4011 ( .A(n3215), .ZN(n3208) );
  INV_X1 U4012 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3332) );
  NAND2_X1 U4013 ( .A1(n4628), .A2(ADDR_REG_2__SCAN_IN), .ZN(n3194) );
  OAI21_X1 U4014 ( .B1(STATE_REG_SCAN_IN), .B2(n3332), .A(n3194), .ZN(n3206)
         );
  OAI211_X1 U4015 ( .C1(n3197), .C2(n3196), .A(n4629), .B(n3195), .ZN(n3204)
         );
  INV_X1 U4016 ( .A(n3198), .ZN(n3202) );
  NAND3_X1 U4017 ( .A1(n3200), .A2(n3199), .A3(n4083), .ZN(n3201) );
  NAND3_X1 U4018 ( .A1(n4587), .A2(n3202), .A3(n3201), .ZN(n3203) );
  NAND2_X1 U4019 ( .A1(n3204), .A2(n3203), .ZN(n3205) );
  AOI211_X1 U4020 ( .C1(n4548), .C2(n4092), .A(n3206), .B(n3205), .ZN(n3207)
         );
  NAND2_X1 U4021 ( .A1(n3208), .A2(n3207), .ZN(U3242) );
  XOR2_X1 U4022 ( .A(REG2_REG_4__SCAN_IN), .B(n3209), .Z(n3217) );
  OAI211_X1 U4023 ( .C1(REG1_REG_4__SCAN_IN), .C2(n3211), .A(n4629), .B(n3210), 
        .ZN(n3213) );
  AND2_X1 U4024 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3780) );
  AOI21_X1 U4025 ( .B1(n4628), .B2(ADDR_REG_4__SCAN_IN), .A(n3780), .ZN(n3212)
         );
  OAI211_X1 U4026 ( .C1(n4635), .C2(n3214), .A(n3213), .B(n3212), .ZN(n3216)
         );
  AOI211_X1 U4027 ( .C1(n4587), .C2(n3217), .A(n3216), .B(n3215), .ZN(n3218)
         );
  INV_X1 U4028 ( .A(n3218), .ZN(U3244) );
  MUX2_X1 U4029 ( .A(REG1_REG_7__SCAN_IN), .B(n4708), .S(n4543), .Z(n3219) );
  XNOR2_X1 U4030 ( .A(n3220), .B(n3219), .ZN(n3229) );
  NOR2_X1 U4031 ( .A1(STATE_REG_SCAN_IN), .A2(n3221), .ZN(n3637) );
  AOI21_X1 U4032 ( .B1(n4628), .B2(ADDR_REG_7__SCAN_IN), .A(n3637), .ZN(n3222)
         );
  OAI21_X1 U4033 ( .B1(n4635), .B2(n3223), .A(n3222), .ZN(n3228) );
  AOI211_X1 U4034 ( .C1(n3226), .C2(n3225), .A(n4622), .B(n3224), .ZN(n3227)
         );
  AOI211_X1 U4035 ( .C1(n4629), .C2(n3229), .A(n3228), .B(n3227), .ZN(n3230)
         );
  INV_X1 U4036 ( .A(n3230), .ZN(U3247) );
  INV_X1 U4037 ( .A(n3231), .ZN(n3234) );
  NAND3_X1 U4038 ( .A1(n3234), .A2(n3233), .A3(n3232), .ZN(n3255) );
  INV_X1 U4039 ( .A(n3255), .ZN(n3248) );
  INV_X1 U4040 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3238) );
  INV_X1 U4041 ( .A(n3885), .ZN(n3823) );
  OAI22_X1 U4042 ( .A1(n3015), .A2(n3823), .B1(n3829), .B2(n3235), .ZN(n3236)
         );
  AOI21_X1 U40430 ( .B1(n3312), .B2(n3887), .A(n3236), .ZN(n3237) );
  OAI21_X1 U4044 ( .B1(n3248), .B2(n3238), .A(n3237), .ZN(U3229) );
  INV_X1 U4045 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3247) );
  INV_X1 U4046 ( .A(n3886), .ZN(n3824) );
  OAI22_X1 U4047 ( .A1(n3239), .A2(n3824), .B1(n3823), .B2(n3017), .ZN(n3240)
         );
  AOI21_X1 U4048 ( .B1(n3241), .B2(n3887), .A(n3240), .ZN(n3246) );
  OAI211_X1 U4049 ( .C1(n3242), .C2(n3244), .A(n3243), .B(n3883), .ZN(n3245)
         );
  OAI211_X1 U4050 ( .C1(n3248), .C2(n3247), .A(n3246), .B(n3245), .ZN(U3219)
         );
  INV_X1 U4051 ( .A(n3249), .ZN(n3250) );
  AOI21_X1 U4052 ( .B1(n3252), .B2(n3251), .A(n3250), .ZN(n3257) );
  AOI22_X1 U4053 ( .A1(n3886), .A2(n4070), .B1(n3885), .B2(n2592), .ZN(n3253)
         );
  OAI21_X1 U4054 ( .B1(n3825), .B2(n3330), .A(n3253), .ZN(n3254) );
  AOI21_X1 U4055 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3255), .A(n3254), .ZN(n3256)
         );
  OAI21_X1 U4056 ( .B1(n3257), .B2(n3829), .A(n3256), .ZN(U3234) );
  XOR2_X1 U4057 ( .A(n3259), .B(n3258), .Z(n3264) );
  OAI22_X1 U4058 ( .A1(n3385), .A2(n3823), .B1(n3824), .B2(n3017), .ZN(n3261)
         );
  MUX2_X1 U4059 ( .A(n3890), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n3260) );
  AOI211_X1 U4060 ( .C1(n3262), .C2(n3887), .A(n3261), .B(n3260), .ZN(n3263)
         );
  OAI21_X1 U4061 ( .B1(n3264), .B2(n3829), .A(n3263), .ZN(U3215) );
  INV_X1 U4062 ( .A(n3266), .ZN(n3911) );
  XNOR2_X1 U4063 ( .A(n3265), .B(n3911), .ZN(n3398) );
  OAI22_X1 U4064 ( .A1(n3017), .A2(n4460), .B1(n3395), .B2(n4459), .ZN(n3269)
         );
  XNOR2_X1 U4065 ( .A(n3267), .B(n3911), .ZN(n3268) );
  OAI22_X1 U4066 ( .A1(n3268), .A2(n4334), .B1(n3385), .B2(n4331), .ZN(n3390)
         );
  AOI211_X1 U4067 ( .C1(n4688), .C2(n3398), .A(n3269), .B(n3390), .ZN(n3274)
         );
  INV_X1 U4068 ( .A(n4467), .ZN(n3348) );
  OR2_X1 U4069 ( .A1(n4678), .A2(n3395), .ZN(n3270) );
  AND2_X1 U4070 ( .A1(n3270), .A2(n3296), .ZN(n3392) );
  AOI22_X1 U4071 ( .A1(n3348), .A2(n3392), .B1(REG1_REG_3__SCAN_IN), .B2(n4710), .ZN(n3271) );
  OAI21_X1 U4072 ( .B1(n3274), .B2(n4710), .A(n3271), .ZN(U3521) );
  NAND2_X1 U4073 ( .A1(n4700), .A2(REG0_REG_3__SCAN_IN), .ZN(n3273) );
  INV_X1 U4074 ( .A(n4531), .ZN(n3346) );
  NAND2_X1 U4075 ( .A1(n3346), .A2(n3392), .ZN(n3272) );
  OAI211_X1 U4076 ( .C1(n3274), .C2(n4700), .A(n3273), .B(n3272), .ZN(U3473)
         );
  OAI21_X1 U4077 ( .B1(n5070), .B2(n3275), .A(n4659), .ZN(n3276) );
  NAND4_X1 U4078 ( .A1(n3279), .A2(n3278), .A3(n3277), .A4(n3276), .ZN(n3280)
         );
  NAND2_X1 U4079 ( .A1(n4648), .A2(n4144), .ZN(n4360) );
  OAI21_X1 U4080 ( .B1(n3310), .B2(n3286), .A(n3329), .ZN(n4673) );
  OR2_X1 U4081 ( .A1(n3056), .A2(n3281), .ZN(n3282) );
  NAND2_X1 U4082 ( .A1(n3283), .A2(n3282), .ZN(n4675) );
  NAND2_X1 U4083 ( .A1(n4072), .A2(n4408), .ZN(n3285) );
  NAND2_X1 U4084 ( .A1(n2574), .A2(n4369), .ZN(n3284) );
  OAI211_X1 U4085 ( .C1(n4459), .C2(n3286), .A(n3285), .B(n3284), .ZN(n3287)
         );
  INV_X1 U4086 ( .A(n3287), .ZN(n3290) );
  XNOR2_X1 U4087 ( .A(n3056), .B(n3931), .ZN(n3288) );
  NAND2_X1 U4088 ( .A1(n3288), .A2(n4367), .ZN(n3289) );
  OAI211_X1 U4089 ( .C1(n4675), .C2(n4312), .A(n3290), .B(n3289), .ZN(n4677)
         );
  MUX2_X1 U4090 ( .A(n4677), .B(REG2_REG_1__SCAN_IN), .S(n4378), .Z(n3291) );
  INV_X1 U4091 ( .A(n3291), .ZN(n3295) );
  INV_X1 U4092 ( .A(n4675), .ZN(n3293) );
  OR2_X1 U4093 ( .A1(n2507), .A2(n4144), .ZN(n3358) );
  INV_X1 U4094 ( .A(n3358), .ZN(n3292) );
  NAND2_X1 U4095 ( .A1(n4648), .A2(n3292), .ZN(n4322) );
  INV_X1 U4096 ( .A(n4322), .ZN(n4653) );
  AOI22_X1 U4097 ( .A1(n3293), .A2(n4653), .B1(REG3_REG_1__SCAN_IN), .B2(n4636), .ZN(n3294) );
  OAI211_X1 U4098 ( .C1(n4385), .C2(n4673), .A(n3295), .B(n3294), .ZN(U3289)
         );
  INV_X1 U4099 ( .A(n3296), .ZN(n3298) );
  OAI211_X1 U4100 ( .C1(n3298), .C2(n3297), .A(n4474), .B(n3344), .ZN(n4683)
         );
  NOR2_X1 U4101 ( .A1(n4683), .A2(n4540), .ZN(n3306) );
  XNOR2_X1 U4102 ( .A(n3299), .B(n3910), .ZN(n3307) );
  XOR2_X1 U4103 ( .A(n3910), .B(n3300), .Z(n3304) );
  AOI22_X1 U4104 ( .A1(n4068), .A2(n4369), .B1(n4406), .B2(n3781), .ZN(n3301)
         );
  OAI21_X1 U4105 ( .B1(n3302), .B2(n4460), .A(n3301), .ZN(n3303) );
  AOI21_X1 U4106 ( .B1(n3304), .B2(n4367), .A(n3303), .ZN(n3305) );
  OAI21_X1 U4107 ( .B1(n3307), .B2(n4312), .A(n3305), .ZN(n4684) );
  AOI211_X1 U4108 ( .C1(n4636), .C2(n3782), .A(n3306), .B(n4684), .ZN(n3309)
         );
  INV_X1 U4109 ( .A(n3307), .ZN(n4686) );
  AOI22_X1 U4110 ( .A1(n4686), .A2(n4653), .B1(REG2_REG_4__SCAN_IN), .B2(n4378), .ZN(n3308) );
  OAI21_X1 U4111 ( .B1(n3309), .B2(n4378), .A(n3308), .ZN(U3286) );
  NAND2_X1 U4112 ( .A1(n4072), .A2(n3310), .ZN(n3933) );
  NAND2_X1 U4113 ( .A1(n3312), .A2(n3311), .ZN(n4669) );
  AOI21_X1 U4114 ( .B1(n4334), .B2(n4312), .A(n4671), .ZN(n3313) );
  AOI21_X1 U4115 ( .B1(n4369), .B2(n4070), .A(n3313), .ZN(n4670) );
  OAI21_X1 U4116 ( .B1(n3314), .B2(n4669), .A(n4670), .ZN(n3315) );
  AOI22_X1 U4117 ( .A1(n3315), .A2(n4648), .B1(REG3_REG_0__SCAN_IN), .B2(n4636), .ZN(n3317) );
  INV_X2 U4118 ( .A(n4648), .ZN(n4378) );
  NAND2_X1 U4119 ( .A1(n4378), .A2(REG2_REG_0__SCAN_IN), .ZN(n3316) );
  OAI211_X1 U4120 ( .C1(n4671), .C2(n4322), .A(n3317), .B(n3316), .ZN(U3290)
         );
  XNOR2_X1 U4121 ( .A(n3318), .B(n3057), .ZN(n3328) );
  NAND2_X1 U4122 ( .A1(n3321), .A2(n3320), .ZN(n3322) );
  NAND2_X1 U4123 ( .A1(n3319), .A2(n3322), .ZN(n4682) );
  INV_X1 U4124 ( .A(n4312), .ZN(n3579) );
  NAND2_X1 U4125 ( .A1(n4682), .A2(n3579), .ZN(n3327) );
  NAND2_X1 U4126 ( .A1(n4070), .A2(n4408), .ZN(n3324) );
  NAND2_X1 U4127 ( .A1(n2592), .A2(n4369), .ZN(n3323) );
  OAI211_X1 U4128 ( .C1(n4459), .C2(n3330), .A(n3324), .B(n3323), .ZN(n3325)
         );
  INV_X1 U4129 ( .A(n3325), .ZN(n3326) );
  OAI211_X1 U4130 ( .C1(n3328), .C2(n4334), .A(n3327), .B(n3326), .ZN(n4680)
         );
  MUX2_X1 U4131 ( .A(n4680), .B(REG2_REG_2__SCAN_IN), .S(n4378), .Z(n3336) );
  NOR2_X1 U4132 ( .A1(n3331), .A2(n3330), .ZN(n4679) );
  NOR3_X1 U4133 ( .A1(n4385), .A2(n4678), .A3(n4679), .ZN(n3335) );
  INV_X1 U4134 ( .A(n4682), .ZN(n3333) );
  OAI22_X1 U4135 ( .A1(n3333), .A2(n4322), .B1(n3332), .B2(n4645), .ZN(n3334)
         );
  OR3_X1 U4136 ( .A1(n3336), .A2(n3335), .A3(n3334), .ZN(U3288) );
  INV_X1 U4137 ( .A(n3338), .ZN(n3944) );
  NAND2_X1 U4138 ( .A1(n3944), .A2(n3961), .ZN(n3922) );
  XOR2_X1 U4139 ( .A(n3337), .B(n3922), .Z(n3387) );
  OAI22_X1 U4140 ( .A1(n3385), .A2(n4460), .B1(n3339), .B2(n4459), .ZN(n3343)
         );
  XOR2_X1 U4141 ( .A(n3922), .B(n3340), .Z(n3342) );
  OAI22_X1 U4142 ( .A1(n3342), .A2(n4334), .B1(n3341), .B2(n4331), .ZN(n3378)
         );
  AOI211_X1 U4143 ( .C1(n3387), .C2(n4688), .A(n3343), .B(n3378), .ZN(n3351)
         );
  AND2_X1 U4144 ( .A1(n3344), .A2(n3749), .ZN(n3345) );
  NOR2_X1 U4145 ( .A1(n2268), .A2(n3345), .ZN(n3382) );
  AOI22_X1 U4146 ( .A1(n3346), .A2(n3382), .B1(REG0_REG_5__SCAN_IN), .B2(n4700), .ZN(n3347) );
  OAI21_X1 U4147 ( .B1(n3351), .B2(n4700), .A(n3347), .ZN(U3477) );
  NAND2_X1 U4148 ( .A1(n4710), .A2(REG1_REG_5__SCAN_IN), .ZN(n3350) );
  NAND2_X1 U4149 ( .A1(n3348), .A2(n3382), .ZN(n3349) );
  OAI211_X1 U4150 ( .C1(n3351), .C2(n4710), .A(n3350), .B(n3349), .ZN(U3523)
         );
  INV_X1 U4151 ( .A(n3920), .ZN(n3948) );
  XNOR2_X1 U4152 ( .A(n3352), .B(n3948), .ZN(n3356) );
  NAND2_X1 U4153 ( .A1(n4067), .A2(n4408), .ZN(n3354) );
  NAND2_X1 U4154 ( .A1(n4065), .A2(n4369), .ZN(n3353) );
  OAI211_X1 U4155 ( .C1(n4459), .C2(n3360), .A(n3354), .B(n3353), .ZN(n3355)
         );
  AOI21_X1 U4156 ( .B1(n3356), .B2(n4367), .A(n3355), .ZN(n4692) );
  XNOR2_X1 U4157 ( .A(n3357), .B(n3948), .ZN(n4689) );
  NAND2_X1 U4158 ( .A1(n4312), .A2(n3358), .ZN(n3359) );
  OAI211_X1 U4159 ( .C1(n2247), .C2(n3360), .A(n4474), .B(n3469), .ZN(n4690)
         );
  NOR2_X1 U4160 ( .A1(n4690), .A2(n4360), .ZN(n3364) );
  INV_X1 U4161 ( .A(n3639), .ZN(n3361) );
  OAI22_X1 U4162 ( .A1(n4648), .A2(n3362), .B1(n3361), .B2(n4645), .ZN(n3363)
         );
  AOI211_X1 U4163 ( .C1(n4689), .C2(n4196), .A(n3364), .B(n3363), .ZN(n3365)
         );
  OAI21_X1 U4164 ( .B1(n4378), .B2(n4692), .A(n3365), .ZN(U3283) );
  AND2_X1 U4165 ( .A1(n3947), .A2(n3959), .ZN(n3902) );
  XNOR2_X1 U4166 ( .A(n3366), .B(n3902), .ZN(n3405) );
  XNOR2_X1 U4167 ( .A(n3367), .B(n3902), .ZN(n3368) );
  AOI22_X1 U4168 ( .A1(n3368), .A2(n4367), .B1(n4369), .B2(n4066), .ZN(n3410)
         );
  AOI22_X1 U4169 ( .A1(n4068), .A2(n4408), .B1(n3861), .B2(n4406), .ZN(n3369)
         );
  OAI211_X1 U4170 ( .C1(n4468), .C2(n3405), .A(n3410), .B(n3369), .ZN(n3376)
         );
  NOR2_X1 U4171 ( .A1(n2268), .A2(n3370), .ZN(n3371) );
  OR2_X1 U4172 ( .A1(n2247), .A2(n3371), .ZN(n3401) );
  INV_X1 U4173 ( .A(REG0_REG_6__SCAN_IN), .ZN(n5010) );
  OAI22_X1 U4174 ( .A1(n3401), .A2(n4531), .B1(n4702), .B2(n5010), .ZN(n3372)
         );
  AOI21_X1 U4175 ( .B1(n3376), .B2(n4702), .A(n3372), .ZN(n3373) );
  INV_X1 U4176 ( .A(n3373), .ZN(U3479) );
  OAI22_X1 U4177 ( .A1(n3401), .A2(n4467), .B1(n4713), .B2(n3374), .ZN(n3375)
         );
  AOI21_X1 U4178 ( .B1(n3376), .B2(n4713), .A(n3375), .ZN(n3377) );
  INV_X1 U4179 ( .A(n3377), .ZN(U3524) );
  INV_X1 U4180 ( .A(n3378), .ZN(n3389) );
  NAND2_X1 U4181 ( .A1(n4648), .A2(n4408), .ZN(n4380) );
  INV_X1 U4182 ( .A(n3750), .ZN(n3379) );
  OAI22_X1 U4183 ( .A1(n4648), .A2(n3380), .B1(n3379), .B2(n4645), .ZN(n3381)
         );
  AOI21_X1 U4184 ( .B1(n3749), .B2(n4382), .A(n3381), .ZN(n3384) );
  NAND2_X1 U4185 ( .A1(n4652), .A2(n3382), .ZN(n3383) );
  OAI211_X1 U4186 ( .C1(n3385), .C2(n4380), .A(n3384), .B(n3383), .ZN(n3386)
         );
  AOI21_X1 U4187 ( .B1(n3387), .B2(n4196), .A(n3386), .ZN(n3388) );
  OAI21_X1 U4188 ( .B1(n3389), .B2(n4378), .A(n3388), .ZN(U3285) );
  INV_X1 U4189 ( .A(n3390), .ZN(n3400) );
  INV_X1 U4190 ( .A(n4382), .ZN(n3396) );
  INV_X1 U4191 ( .A(n4380), .ZN(n3494) );
  INV_X1 U4192 ( .A(REG2_REG_3__SCAN_IN), .ZN(n4095) );
  OAI22_X1 U4193 ( .A1(n4648), .A2(n4095), .B1(REG3_REG_3__SCAN_IN), .B2(n4645), .ZN(n3391) );
  AOI21_X1 U4194 ( .B1(n3494), .B2(n2574), .A(n3391), .ZN(n3394) );
  NAND2_X1 U4195 ( .A1(n4652), .A2(n3392), .ZN(n3393) );
  OAI211_X1 U4196 ( .C1(n3396), .C2(n3395), .A(n3394), .B(n3393), .ZN(n3397)
         );
  AOI21_X1 U4197 ( .B1(n3398), .B2(n4196), .A(n3397), .ZN(n3399) );
  OAI21_X1 U4198 ( .B1(n3400), .B2(n4378), .A(n3399), .ZN(U3287) );
  INV_X1 U4199 ( .A(n3401), .ZN(n3408) );
  AOI22_X1 U4200 ( .A1(n4378), .A2(REG2_REG_6__SCAN_IN), .B1(n3862), .B2(n4636), .ZN(n3403) );
  NAND2_X1 U4201 ( .A1(n4382), .A2(n3861), .ZN(n3402) );
  OAI211_X1 U4202 ( .C1(n3404), .C2(n4380), .A(n3403), .B(n3402), .ZN(n3407)
         );
  NOR2_X1 U4203 ( .A1(n3405), .A2(n4388), .ZN(n3406) );
  AOI211_X1 U4204 ( .C1(n3408), .C2(n4652), .A(n3407), .B(n3406), .ZN(n3409)
         );
  OAI21_X1 U4205 ( .B1(n4378), .B2(n3410), .A(n3409), .ZN(U3284) );
  INV_X1 U4206 ( .A(n3969), .ZN(n3411) );
  NAND2_X1 U4207 ( .A1(n3411), .A2(n3952), .ZN(n3919) );
  XOR2_X1 U4208 ( .A(n3412), .B(n3919), .Z(n3414) );
  OAI22_X1 U4209 ( .A1(n3414), .A2(n4334), .B1(n3413), .B2(n4331), .ZN(n3461)
         );
  INV_X1 U4210 ( .A(n3461), .ZN(n3424) );
  XNOR2_X1 U4211 ( .A(n3415), .B(n3919), .ZN(n3463) );
  AND2_X1 U4212 ( .A1(n3470), .A2(n3790), .ZN(n3416) );
  OR2_X1 U4213 ( .A1(n3416), .A2(n3531), .ZN(n3468) );
  INV_X1 U4214 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3417) );
  OAI22_X1 U4215 ( .A1(n3418), .A2(n4645), .B1(n3417), .B2(n4648), .ZN(n3419)
         );
  AOI21_X1 U4216 ( .B1(n4382), .B2(n3790), .A(n3419), .ZN(n3421) );
  OR2_X1 U4217 ( .A1(n4380), .A2(n3460), .ZN(n3420) );
  OAI211_X1 U4218 ( .C1(n3468), .C2(n4385), .A(n3421), .B(n3420), .ZN(n3422)
         );
  AOI21_X1 U4219 ( .B1(n3463), .B2(n4196), .A(n3422), .ZN(n3423) );
  OAI21_X1 U4220 ( .B1(n3424), .B2(n4378), .A(n3423), .ZN(U3281) );
  INV_X1 U4221 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4711) );
  AOI22_X1 U4222 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3443), .B1(n4667), .B2(
        n4711), .ZN(n4577) );
  NAND2_X1 U4223 ( .A1(n4553), .A2(REG1_REG_9__SCAN_IN), .ZN(n3430) );
  INV_X1 U4224 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3425) );
  MUX2_X1 U4225 ( .A(n3425), .B(REG1_REG_9__SCAN_IN), .S(n4553), .Z(n3426) );
  INV_X1 U4226 ( .A(n3426), .ZN(n4558) );
  INV_X1 U4227 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3427) );
  OAI22_X1 U4228 ( .A1(n3429), .A2(n3444), .B1(n3428), .B2(n3427), .ZN(n4559)
         );
  NAND2_X1 U4229 ( .A1(n4558), .A2(n4559), .ZN(n4557) );
  NAND2_X1 U4230 ( .A1(n3430), .A2(n4557), .ZN(n3431) );
  NAND2_X1 U4231 ( .A1(n3448), .A2(n3431), .ZN(n3432) );
  INV_X1 U4232 ( .A(n3448), .ZN(n4668) );
  XNOR2_X1 U4233 ( .A(n3431), .B(n4668), .ZN(n4572) );
  NAND2_X1 U4234 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4572), .ZN(n4571) );
  NAND2_X1 U4235 ( .A1(n3432), .A2(n4571), .ZN(n4576) );
  NAND2_X1 U4236 ( .A1(n4577), .A2(n4576), .ZN(n4575) );
  OAI21_X1 U4237 ( .B1(n4667), .B2(n4711), .A(n4575), .ZN(n3433) );
  NAND2_X1 U4238 ( .A1(n3452), .A2(n3433), .ZN(n3434) );
  INV_X1 U4239 ( .A(n3452), .ZN(n4665) );
  XNOR2_X1 U4240 ( .A(n3433), .B(n4665), .ZN(n4593) );
  NAND2_X1 U4241 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4593), .ZN(n4592) );
  NAND2_X1 U4242 ( .A1(n3434), .A2(n4592), .ZN(n3436) );
  INV_X1 U4243 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3591) );
  NOR2_X1 U4244 ( .A1(n3440), .A2(n3591), .ZN(n4102) );
  AOI21_X1 U4245 ( .B1(n3591), .B2(n3440), .A(n4102), .ZN(n3435) );
  NAND2_X1 U4246 ( .A1(n3435), .A2(n3436), .ZN(n4103) );
  OAI211_X1 U4247 ( .C1(n3436), .C2(n3435), .A(n4629), .B(n4103), .ZN(n3439)
         );
  INV_X1 U4248 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3437) );
  NOR2_X1 U4249 ( .A1(STATE_REG_SCAN_IN), .A2(n3437), .ZN(n3812) );
  AOI21_X1 U4250 ( .B1(n4628), .B2(ADDR_REG_13__SCAN_IN), .A(n3812), .ZN(n3438) );
  OAI211_X1 U4251 ( .C1(n4635), .C2(n3440), .A(n3439), .B(n3438), .ZN(n3458)
         );
  INV_X1 U4252 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3441) );
  NOR2_X1 U4253 ( .A1(n3440), .A2(n3441), .ZN(n4117) );
  AOI21_X1 U4254 ( .B1(n3441), .B2(n3440), .A(n4117), .ZN(n3456) );
  NAND2_X1 U4255 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3443), .ZN(n3451) );
  INV_X1 U4256 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3442) );
  AOI22_X1 U4257 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3443), .B1(n4667), .B2(
        n3442), .ZN(n4580) );
  NAND2_X1 U4258 ( .A1(n4553), .A2(REG2_REG_9__SCAN_IN), .ZN(n3447) );
  MUX2_X1 U4259 ( .A(REG2_REG_9__SCAN_IN), .B(n3417), .S(n4553), .Z(n4555) );
  INV_X1 U4260 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4647) );
  OAI22_X1 U4261 ( .A1(n3446), .A2(n4647), .B1(n3445), .B2(n3444), .ZN(n4556)
         );
  NAND2_X1 U4262 ( .A1(n4555), .A2(n4556), .ZN(n4554) );
  NAND2_X1 U4263 ( .A1(n3447), .A2(n4554), .ZN(n3449) );
  NAND2_X1 U4264 ( .A1(n3448), .A2(n3449), .ZN(n3450) );
  XNOR2_X1 U4265 ( .A(n3449), .B(n4668), .ZN(n4567) );
  NAND2_X1 U4266 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4567), .ZN(n4566) );
  NAND2_X1 U4267 ( .A1(n3450), .A2(n4566), .ZN(n4579) );
  NAND2_X1 U4268 ( .A1(n4580), .A2(n4579), .ZN(n4578) );
  NAND2_X1 U4269 ( .A1(n3452), .A2(n3453), .ZN(n3454) );
  OAI21_X1 U4270 ( .B1(n3456), .B2(n4118), .A(n4587), .ZN(n3455) );
  AOI21_X1 U4271 ( .B1(n3456), .B2(n4118), .A(n3455), .ZN(n3457) );
  OR2_X1 U4272 ( .A1(n3458), .A2(n3457), .ZN(U3253) );
  INV_X1 U4273 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3464) );
  OAI22_X1 U4274 ( .A1(n3460), .A2(n4460), .B1(n3459), .B2(n4459), .ZN(n3462)
         );
  AOI211_X1 U4275 ( .C1(n4688), .C2(n3463), .A(n3462), .B(n3461), .ZN(n3466)
         );
  MUX2_X1 U4276 ( .A(n3464), .B(n3466), .S(n4702), .Z(n3465) );
  OAI21_X1 U4277 ( .B1(n3468), .B2(n4531), .A(n3465), .ZN(U3485) );
  MUX2_X1 U4278 ( .A(n3425), .B(n3466), .S(n4713), .Z(n3467) );
  OAI21_X1 U4279 ( .B1(n4467), .B2(n3468), .A(n3467), .ZN(U3527) );
  INV_X1 U4280 ( .A(n3469), .ZN(n3471) );
  OAI21_X1 U4281 ( .B1(n3471), .B2(n3474), .A(n3470), .ZN(n4650) );
  INV_X1 U4282 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3481) );
  NAND2_X1 U4283 ( .A1(n3953), .A2(n3950), .ZN(n3917) );
  XOR2_X1 U4284 ( .A(n3917), .B(n3472), .Z(n4654) );
  XOR2_X1 U4285 ( .A(n3473), .B(n3917), .Z(n3478) );
  OAI22_X1 U4286 ( .A1(n3475), .A2(n4460), .B1(n3474), .B2(n4459), .ZN(n3476)
         );
  AOI21_X1 U4287 ( .B1(n4369), .B2(n4064), .A(n3476), .ZN(n3477) );
  OAI21_X1 U4288 ( .B1(n3478), .B2(n4334), .A(n3477), .ZN(n3479) );
  AOI21_X1 U4289 ( .B1(n3579), .B2(n4654), .A(n3479), .ZN(n4657) );
  INV_X1 U4290 ( .A(n4657), .ZN(n3480) );
  AOI21_X1 U4291 ( .B1(n4699), .B2(n4654), .A(n3480), .ZN(n3483) );
  MUX2_X1 U4292 ( .A(n3481), .B(n3483), .S(n4702), .Z(n3482) );
  OAI21_X1 U4293 ( .B1(n4650), .B2(n4531), .A(n3482), .ZN(U3483) );
  MUX2_X1 U4294 ( .A(n3427), .B(n3483), .S(n4713), .Z(n3484) );
  OAI21_X1 U4295 ( .B1(n4650), .B2(n4467), .A(n3484), .ZN(U3526) );
  NAND2_X1 U4296 ( .A1(n3515), .A2(n3513), .ZN(n3918) );
  INV_X1 U4297 ( .A(n3485), .ZN(n3486) );
  AOI21_X1 U4298 ( .B1(n3500), .B2(n3487), .A(n3486), .ZN(n3516) );
  XOR2_X1 U4299 ( .A(n3918), .B(n3516), .Z(n3488) );
  OAI22_X1 U4300 ( .A1(n3488), .A2(n4334), .B1(n3577), .B2(n4331), .ZN(n3548)
         );
  INV_X1 U4301 ( .A(n3548), .ZN(n3499) );
  XNOR2_X1 U4302 ( .A(n3489), .B(n3918), .ZN(n3550) );
  NAND2_X1 U4303 ( .A1(n3507), .A2(n3720), .ZN(n3490) );
  NAND2_X1 U4304 ( .A1(n3523), .A2(n3490), .ZN(n3556) );
  INV_X1 U4305 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3492) );
  INV_X1 U4306 ( .A(n3721), .ZN(n3491) );
  OAI22_X1 U4307 ( .A1(n4648), .A2(n3492), .B1(n3491), .B2(n4645), .ZN(n3493)
         );
  AOI21_X1 U4308 ( .B1(n3494), .B2(n4062), .A(n3493), .ZN(n3496) );
  NAND2_X1 U4309 ( .A1(n4382), .A2(n3720), .ZN(n3495) );
  OAI211_X1 U4310 ( .C1(n3556), .C2(n4385), .A(n3496), .B(n3495), .ZN(n3497)
         );
  AOI21_X1 U4311 ( .B1(n3550), .B2(n4196), .A(n3497), .ZN(n3498) );
  OAI21_X1 U4312 ( .B1(n3499), .B2(n4378), .A(n3498), .ZN(U3278) );
  XNOR2_X1 U4313 ( .A(n3500), .B(n3921), .ZN(n3506) );
  XNOR2_X1 U4314 ( .A(n3501), .B(n3921), .ZN(n4698) );
  NAND2_X1 U4315 ( .A1(n4698), .A2(n3579), .ZN(n3505) );
  OAI22_X1 U4316 ( .A1(n3502), .A2(n4331), .B1(n4459), .B2(n3508), .ZN(n3503)
         );
  AOI21_X1 U4317 ( .B1(n4408), .B2(n4063), .A(n3503), .ZN(n3504) );
  OAI211_X1 U4318 ( .C1(n4334), .C2(n3506), .A(n3505), .B(n3504), .ZN(n4696)
         );
  INV_X1 U4319 ( .A(n4696), .ZN(n3512) );
  OAI21_X1 U4320 ( .B1(n3529), .B2(n3508), .A(n3507), .ZN(n4695) );
  AOI22_X1 U4321 ( .A1(n4378), .A2(REG2_REG_11__SCAN_IN), .B1(n3838), .B2(
        n4636), .ZN(n3509) );
  OAI21_X1 U4322 ( .B1(n4695), .B2(n4385), .A(n3509), .ZN(n3510) );
  AOI21_X1 U4323 ( .B1(n4698), .B2(n4653), .A(n3510), .ZN(n3511) );
  OAI21_X1 U4324 ( .B1(n3512), .B2(n4378), .A(n3511), .ZN(U3279) );
  INV_X1 U4325 ( .A(n3513), .ZN(n3514) );
  AOI21_X1 U4326 ( .B1(n3516), .B2(n3515), .A(n3514), .ZN(n3517) );
  XNOR2_X1 U4327 ( .A(n4060), .B(n3518), .ZN(n3928) );
  XNOR2_X1 U4328 ( .A(n3517), .B(n3928), .ZN(n3521) );
  OAI22_X1 U4329 ( .A1(n3595), .A2(n4331), .B1(n4459), .B2(n3518), .ZN(n3519)
         );
  AOI21_X1 U4330 ( .B1(n4408), .B2(n4061), .A(n3519), .ZN(n3520) );
  OAI21_X1 U4331 ( .B1(n3521), .B2(n4334), .A(n3520), .ZN(n3586) );
  INV_X1 U4332 ( .A(n3586), .ZN(n3528) );
  XOR2_X1 U4333 ( .A(n3928), .B(n3522), .Z(n3587) );
  AND2_X1 U4334 ( .A1(n3523), .A2(n3813), .ZN(n3524) );
  OR2_X1 U4335 ( .A1(n3524), .A2(n2238), .ZN(n3593) );
  AOI22_X1 U4336 ( .A1(n4378), .A2(REG2_REG_13__SCAN_IN), .B1(n3814), .B2(
        n4636), .ZN(n3525) );
  OAI21_X1 U4337 ( .B1(n3593), .B2(n4385), .A(n3525), .ZN(n3526) );
  AOI21_X1 U4338 ( .B1(n3587), .B2(n4196), .A(n3526), .ZN(n3527) );
  OAI21_X1 U4339 ( .B1(n4378), .B2(n3528), .A(n3527), .ZN(U3277) );
  INV_X1 U4340 ( .A(n3529), .ZN(n3530) );
  OAI21_X1 U4341 ( .B1(n3531), .B2(n3534), .A(n3530), .ZN(n4638) );
  INV_X1 U4342 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3541) );
  AND2_X1 U4343 ( .A1(n3970), .A2(n3972), .ZN(n3903) );
  XNOR2_X1 U4344 ( .A(n3532), .B(n3903), .ZN(n4640) );
  XOR2_X1 U4345 ( .A(n3533), .B(n3903), .Z(n3538) );
  OAI22_X1 U4346 ( .A1(n3535), .A2(n4460), .B1(n3534), .B2(n4459), .ZN(n3536)
         );
  AOI21_X1 U4347 ( .B1(n4369), .B2(n4062), .A(n3536), .ZN(n3537) );
  OAI21_X1 U4348 ( .B1(n3538), .B2(n4334), .A(n3537), .ZN(n3539) );
  AOI21_X1 U4349 ( .B1(n3579), .B2(n4640), .A(n3539), .ZN(n4643) );
  INV_X1 U4350 ( .A(n4643), .ZN(n3540) );
  AOI21_X1 U4351 ( .B1(n4699), .B2(n4640), .A(n3540), .ZN(n3543) );
  MUX2_X1 U4352 ( .A(n3541), .B(n3543), .S(n4702), .Z(n3542) );
  OAI21_X1 U4353 ( .B1(n4638), .B2(n4531), .A(n3542), .ZN(U3487) );
  INV_X1 U4354 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3544) );
  MUX2_X1 U4355 ( .A(n3544), .B(n3543), .S(n4713), .Z(n3545) );
  OAI21_X1 U4356 ( .B1(n4638), .B2(n4467), .A(n3545), .ZN(U3528) );
  INV_X1 U4357 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3551) );
  OAI22_X1 U4358 ( .A1(n3547), .A2(n4460), .B1(n3546), .B2(n4459), .ZN(n3549)
         );
  AOI211_X1 U4359 ( .C1(n4688), .C2(n3550), .A(n3549), .B(n3548), .ZN(n3553)
         );
  MUX2_X1 U4360 ( .A(n3551), .B(n3553), .S(n4713), .Z(n3552) );
  OAI21_X1 U4361 ( .B1(n3556), .B2(n4467), .A(n3552), .ZN(U3530) );
  INV_X1 U4362 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3554) );
  MUX2_X1 U4363 ( .A(n3554), .B(n3553), .S(n4702), .Z(n3555) );
  OAI21_X1 U4364 ( .B1(n3556), .B2(n4531), .A(n3555), .ZN(U3491) );
  XNOR2_X1 U4365 ( .A(n3557), .B(n3905), .ZN(n3598) );
  INV_X1 U4366 ( .A(n3598), .ZN(n3569) );
  NAND2_X1 U4367 ( .A1(n3572), .A2(n3977), .ZN(n3559) );
  INV_X1 U4368 ( .A(n3905), .ZN(n3558) );
  XNOR2_X1 U4369 ( .A(n3559), .B(n3558), .ZN(n3560) );
  NAND2_X1 U4370 ( .A1(n3560), .A2(n4367), .ZN(n3562) );
  NAND2_X1 U4371 ( .A1(n4057), .A2(n4369), .ZN(n3561) );
  NAND2_X1 U4372 ( .A1(n3562), .A2(n3561), .ZN(n3597) );
  INV_X1 U4373 ( .A(n4476), .ZN(n3563) );
  OAI21_X1 U4374 ( .B1(n3563), .B2(n3594), .A(n3607), .ZN(n3604) );
  AOI22_X1 U4375 ( .A1(n4378), .A2(REG2_REG_15__SCAN_IN), .B1(n3889), .B2(
        n4636), .ZN(n3564) );
  OAI21_X1 U4376 ( .B1(n3595), .B2(n4380), .A(n3564), .ZN(n3565) );
  AOI21_X1 U4377 ( .B1(n3888), .B2(n4382), .A(n3565), .ZN(n3566) );
  OAI21_X1 U4378 ( .B1(n3604), .B2(n4385), .A(n3566), .ZN(n3567) );
  AOI21_X1 U4379 ( .B1(n3597), .B2(n4648), .A(n3567), .ZN(n3568) );
  OAI21_X1 U4380 ( .B1(n3569), .B2(n4388), .A(n3568), .ZN(U3275) );
  OAI21_X1 U4381 ( .B1(n3571), .B2(n3906), .A(n3570), .ZN(n3580) );
  OAI21_X1 U4382 ( .B1(n3573), .B2(n4011), .A(n3572), .ZN(n3574) );
  NAND2_X1 U4383 ( .A1(n3574), .A2(n4367), .ZN(n3576) );
  AOI22_X1 U4384 ( .A1(n4058), .A2(n4369), .B1(n4406), .B2(n3656), .ZN(n3575)
         );
  OAI211_X1 U4385 ( .C1(n3577), .C2(n4460), .A(n3576), .B(n3575), .ZN(n3578)
         );
  AOI21_X1 U4386 ( .B1(n3580), .B2(n3579), .A(n3578), .ZN(n4478) );
  INV_X1 U4387 ( .A(n3580), .ZN(n4479) );
  AOI22_X1 U4388 ( .A1(n4378), .A2(REG2_REG_14__SCAN_IN), .B1(n3657), .B2(
        n4636), .ZN(n3583) );
  OR2_X1 U4389 ( .A1(n2238), .A2(n3581), .ZN(n4475) );
  NAND3_X1 U4390 ( .A1(n4476), .A2(n4475), .A3(n4652), .ZN(n3582) );
  OAI211_X1 U4391 ( .C1(n4479), .C2(n4322), .A(n3583), .B(n3582), .ZN(n3584)
         );
  INV_X1 U4392 ( .A(n3584), .ZN(n3585) );
  OAI21_X1 U4393 ( .B1(n4378), .B2(n4478), .A(n3585), .ZN(U3276) );
  INV_X1 U4394 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3588) );
  AOI21_X1 U4395 ( .B1(n3587), .B2(n4688), .A(n3586), .ZN(n3590) );
  MUX2_X1 U4396 ( .A(n3588), .B(n3590), .S(n4702), .Z(n3589) );
  OAI21_X1 U4397 ( .B1(n3593), .B2(n4531), .A(n3589), .ZN(U3493) );
  MUX2_X1 U4398 ( .A(n3591), .B(n3590), .S(n4713), .Z(n3592) );
  OAI21_X1 U4399 ( .B1(n4467), .B2(n3593), .A(n3592), .ZN(U3531) );
  INV_X1 U4400 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3599) );
  OAI22_X1 U4401 ( .A1(n3595), .A2(n4460), .B1(n3594), .B2(n4459), .ZN(n3596)
         );
  AOI211_X1 U4402 ( .C1(n3598), .C2(n4688), .A(n3597), .B(n3596), .ZN(n3601)
         );
  MUX2_X1 U4403 ( .A(n3599), .B(n3601), .S(n4702), .Z(n3600) );
  OAI21_X1 U4404 ( .B1(n3604), .B2(n4531), .A(n3600), .ZN(U3497) );
  INV_X1 U4405 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3602) );
  MUX2_X1 U4406 ( .A(n3602), .B(n3601), .S(n4713), .Z(n3603) );
  OAI21_X1 U4407 ( .B1(n4467), .B2(n3604), .A(n3603), .ZN(U3533) );
  OAI21_X1 U4408 ( .B1(n3606), .B2(n3613), .A(n3605), .ZN(n4469) );
  NAND2_X1 U4409 ( .A1(n3607), .A2(n3739), .ZN(n3608) );
  NAND2_X1 U4410 ( .A1(n4373), .A2(n3608), .ZN(n4534) );
  INV_X1 U4411 ( .A(n4534), .ZN(n3612) );
  INV_X1 U4412 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3610) );
  INV_X1 U4413 ( .A(n3740), .ZN(n3609) );
  OAI22_X1 U4414 ( .A1(n4648), .A2(n3610), .B1(n3609), .B2(n4645), .ZN(n3611)
         );
  AOI21_X1 U4415 ( .B1(n3612), .B2(n4652), .A(n3611), .ZN(n3621) );
  XNOR2_X1 U4416 ( .A(n3614), .B(n3613), .ZN(n3619) );
  NAND2_X1 U4417 ( .A1(n4058), .A2(n4408), .ZN(n3616) );
  NAND2_X1 U4418 ( .A1(n4056), .A2(n4369), .ZN(n3615) );
  OAI211_X1 U4419 ( .C1(n4459), .C2(n3617), .A(n3616), .B(n3615), .ZN(n3618)
         );
  AOI21_X1 U4420 ( .B1(n3619), .B2(n4367), .A(n3618), .ZN(n4470) );
  OR2_X1 U4421 ( .A1(n4470), .A2(n4378), .ZN(n3620) );
  OAI211_X1 U4422 ( .C1(n4469), .C2(n4388), .A(n3621), .B(n3620), .ZN(U3274)
         );
  INV_X1 U4423 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3623) );
  OAI22_X1 U4424 ( .A1(n3624), .A2(n4380), .B1(n3623), .B2(n4648), .ZN(n3625)
         );
  AOI21_X1 U4425 ( .B1(n4000), .B2(n4382), .A(n3625), .ZN(n3631) );
  OAI22_X1 U4426 ( .A1(n3627), .A2(n4385), .B1(n3626), .B2(n4645), .ZN(n3628)
         );
  OAI21_X1 U4427 ( .B1(n3629), .B2(n3628), .A(n4648), .ZN(n3630) );
  OAI211_X1 U4428 ( .C1(n3622), .C2(n4388), .A(n3631), .B(n3630), .ZN(U3354)
         );
  INV_X1 U4429 ( .A(IR_REG_30__SCAN_IN), .ZN(n3632) );
  NAND3_X1 U4430 ( .A1(n3632), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3633) );
  INV_X1 U4431 ( .A(DATAI_31_), .ZN(n4827) );
  OAI22_X1 U4432 ( .A1(n2471), .A2(n3633), .B1(STATE_REG_SCAN_IN), .B2(n4827), 
        .ZN(U3321) );
  XOR2_X1 U4433 ( .A(n3634), .B(n3635), .Z(n3636) );
  NAND2_X1 U4434 ( .A1(n3636), .A2(n3883), .ZN(n3643) );
  AOI21_X1 U4435 ( .B1(n3886), .B2(n4067), .A(n3637), .ZN(n3642) );
  AOI22_X1 U4436 ( .A1(n3638), .A2(n3887), .B1(n3885), .B2(n4065), .ZN(n3641)
         );
  NAND2_X1 U4437 ( .A1(n3890), .A2(n3639), .ZN(n3640) );
  NAND4_X1 U4438 ( .A1(n3643), .A2(n3642), .A3(n3641), .A4(n3640), .ZN(U3210)
         );
  XNOR2_X1 U4439 ( .A(n3644), .B(n2257), .ZN(n3645) );
  NAND2_X1 U4440 ( .A1(n3645), .A2(n3883), .ZN(n3649) );
  AOI22_X1 U4441 ( .A1(n4179), .A2(n3885), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3648) );
  AOI22_X1 U4442 ( .A1(n4407), .A2(n3887), .B1(n3886), .B2(n4409), .ZN(n3647)
         );
  NAND2_X1 U4443 ( .A1(n3890), .A2(n4173), .ZN(n3646) );
  NAND4_X1 U4444 ( .A1(n3649), .A2(n3648), .A3(n3647), .A4(n3646), .ZN(U3211)
         );
  INV_X1 U4445 ( .A(n3650), .ZN(n3652) );
  NAND2_X1 U4446 ( .A1(n3652), .A2(n3651), .ZN(n3653) );
  XNOR2_X1 U4447 ( .A(n3654), .B(n3653), .ZN(n3655) );
  NAND2_X1 U4448 ( .A1(n3655), .A2(n3883), .ZN(n3661) );
  AND2_X1 U4449 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4600) );
  AOI21_X1 U4450 ( .B1(n3886), .B2(n4060), .A(n4600), .ZN(n3660) );
  AOI22_X1 U4451 ( .A1(n3656), .A2(n3887), .B1(n3885), .B2(n4058), .ZN(n3659)
         );
  NAND2_X1 U4452 ( .A1(n3890), .A2(n3657), .ZN(n3658) );
  NAND4_X1 U4453 ( .A1(n3661), .A2(n3660), .A3(n3659), .A4(n3658), .ZN(U3212)
         );
  OAI21_X1 U4454 ( .B1(n3819), .B2(n3663), .A(n3662), .ZN(n3664) );
  NAND3_X1 U4455 ( .A1(n2253), .A2(n3883), .A3(n3664), .ZN(n3668) );
  AOI22_X1 U4456 ( .A1(n3885), .A2(n4212), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3667) );
  AOI22_X1 U4457 ( .A1(n4260), .A2(n3887), .B1(n3886), .B2(n4257), .ZN(n3666)
         );
  NAND2_X1 U4458 ( .A1(n3890), .A2(n4263), .ZN(n3665) );
  NAND4_X1 U4459 ( .A1(n3668), .A2(n3667), .A3(n3666), .A4(n3665), .ZN(U3213)
         );
  AOI21_X1 U4460 ( .B1(n3669), .B2(n3670), .A(n3829), .ZN(n3672) );
  NAND2_X1 U4461 ( .A1(n3672), .A2(n3671), .ZN(n3678) );
  NAND2_X1 U4462 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4568) );
  INV_X1 U4463 ( .A(n4568), .ZN(n3673) );
  AOI21_X1 U4464 ( .B1(n3886), .B2(n4064), .A(n3673), .ZN(n3677) );
  AOI22_X1 U4465 ( .A1(n3674), .A2(n3887), .B1(n3885), .B2(n4062), .ZN(n3676)
         );
  NAND2_X1 U4466 ( .A1(n3890), .A2(n4637), .ZN(n3675) );
  NAND4_X1 U4467 ( .A1(n3678), .A2(n3677), .A3(n3676), .A4(n3675), .ZN(U3214)
         );
  XNOR2_X1 U4468 ( .A(n3680), .B(n3679), .ZN(n3681) );
  NAND2_X1 U4469 ( .A1(n3681), .A2(n3883), .ZN(n3687) );
  NAND2_X1 U4470 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4143) );
  INV_X1 U4471 ( .A(n4143), .ZN(n3682) );
  AOI21_X1 U4472 ( .B1(n3885), .B2(n4055), .A(n3682), .ZN(n3686) );
  AOI22_X1 U4473 ( .A1(n3683), .A2(n3887), .B1(n3886), .B2(n4370), .ZN(n3685)
         );
  NAND2_X1 U4474 ( .A1(n3890), .A2(n4339), .ZN(n3684) );
  NAND4_X1 U4475 ( .A1(n3687), .A2(n3686), .A3(n3685), .A4(n3684), .ZN(U3216)
         );
  INV_X1 U4476 ( .A(n3689), .ZN(n3691) );
  NAND2_X1 U4477 ( .A1(n3691), .A2(n3690), .ZN(n3692) );
  XNOR2_X1 U4478 ( .A(n3688), .B(n3692), .ZN(n3693) );
  NAND2_X1 U4479 ( .A1(n3693), .A2(n3883), .ZN(n3700) );
  INV_X1 U4480 ( .A(n3694), .ZN(n3695) );
  AOI21_X1 U4481 ( .B1(n3886), .B2(n4066), .A(n3695), .ZN(n3699) );
  AOI22_X1 U4482 ( .A1(n3696), .A2(n3887), .B1(n3885), .B2(n4064), .ZN(n3698)
         );
  NAND2_X1 U4483 ( .A1(n3890), .A2(n4644), .ZN(n3697) );
  NAND4_X1 U4484 ( .A1(n3700), .A2(n3699), .A3(n3698), .A4(n3697), .ZN(U3218)
         );
  AOI21_X1 U4485 ( .B1(n3800), .B2(n3797), .A(n3796), .ZN(n3705) );
  XOR2_X1 U4486 ( .A(n3703), .B(n3702), .Z(n3704) );
  XNOR2_X1 U4487 ( .A(n3705), .B(n3704), .ZN(n3706) );
  NAND2_X1 U4488 ( .A1(n3706), .A2(n3883), .ZN(n3710) );
  AOI22_X1 U4489 ( .A1(n3885), .A2(n4257), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3709) );
  AOI22_X1 U4490 ( .A1(n4296), .A2(n3887), .B1(n3886), .B2(n4055), .ZN(n3708)
         );
  NAND2_X1 U4491 ( .A1(n3890), .A2(n4293), .ZN(n3707) );
  NAND4_X1 U4492 ( .A1(n3710), .A2(n3709), .A3(n3708), .A4(n3707), .ZN(U3220)
         );
  INV_X1 U4493 ( .A(n3831), .ZN(n3711) );
  NOR2_X1 U4494 ( .A1(n3834), .A2(n3711), .ZN(n3713) );
  OAI22_X1 U4495 ( .A1(n3713), .A2(n3832), .B1(n3712), .B2(n3831), .ZN(n3717)
         );
  NAND2_X1 U4496 ( .A1(n3715), .A2(n3714), .ZN(n3716) );
  XNOR2_X1 U4497 ( .A(n3717), .B(n3716), .ZN(n3718) );
  NAND2_X1 U4498 ( .A1(n3718), .A2(n3883), .ZN(n3725) );
  NAND2_X1 U4499 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4589) );
  INV_X1 U4500 ( .A(n4589), .ZN(n3719) );
  AOI21_X1 U4501 ( .B1(n3886), .B2(n4062), .A(n3719), .ZN(n3724) );
  AOI22_X1 U4502 ( .A1(n3720), .A2(n3887), .B1(n3885), .B2(n4060), .ZN(n3723)
         );
  NAND2_X1 U4503 ( .A1(n3890), .A2(n3721), .ZN(n3722) );
  NAND4_X1 U4504 ( .A1(n3725), .A2(n3724), .A3(n3723), .A4(n3722), .ZN(U3221)
         );
  INV_X1 U4505 ( .A(n3726), .ZN(n3728) );
  NAND2_X1 U4506 ( .A1(n3728), .A2(n3727), .ZN(n3729) );
  XNOR2_X1 U4507 ( .A(n3730), .B(n3729), .ZN(n3731) );
  NAND2_X1 U4508 ( .A1(n3731), .A2(n3883), .ZN(n3735) );
  AOI22_X1 U4509 ( .A1(n3885), .A2(n4409), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3734) );
  AOI22_X1 U4510 ( .A1(n4211), .A2(n3887), .B1(n3886), .B2(n4212), .ZN(n3733)
         );
  NAND2_X1 U4511 ( .A1(n3890), .A2(n4221), .ZN(n3732) );
  NAND4_X1 U4512 ( .A1(n3735), .A2(n3734), .A3(n3733), .A4(n3732), .ZN(U3222)
         );
  OAI21_X1 U4513 ( .B1(n3878), .B2(n3881), .A(n3879), .ZN(n3736) );
  XOR2_X1 U4514 ( .A(n3737), .B(n3736), .Z(n3738) );
  NAND2_X1 U4515 ( .A1(n3738), .A2(n3883), .ZN(n3744) );
  NOR2_X1 U4516 ( .A1(STATE_REG_SCAN_IN), .A2(n5073), .ZN(n4617) );
  AOI21_X1 U4517 ( .B1(n3885), .B2(n4056), .A(n4617), .ZN(n3743) );
  AOI22_X1 U4518 ( .A1(n3739), .A2(n3887), .B1(n3886), .B2(n4058), .ZN(n3742)
         );
  NAND2_X1 U4519 ( .A1(n3890), .A2(n3740), .ZN(n3741) );
  NAND4_X1 U4520 ( .A1(n3744), .A2(n3743), .A3(n3742), .A4(n3741), .ZN(U3223)
         );
  OAI211_X1 U4521 ( .C1(n3747), .C2(n3746), .A(n3745), .B(n3883), .ZN(n3754)
         );
  AOI21_X1 U4522 ( .B1(n3886), .B2(n4069), .A(n3748), .ZN(n3753) );
  AOI22_X1 U4523 ( .A1(n3749), .A2(n3887), .B1(n3885), .B2(n4067), .ZN(n3752)
         );
  NAND2_X1 U4524 ( .A1(n3890), .A2(n3750), .ZN(n3751) );
  NAND4_X1 U4525 ( .A1(n3754), .A2(n3753), .A3(n3752), .A4(n3751), .ZN(U3224)
         );
  INV_X1 U4526 ( .A(n3755), .ZN(n3757) );
  NAND2_X1 U4527 ( .A1(n3757), .A2(n3756), .ZN(n3758) );
  XNOR2_X1 U4528 ( .A(n3759), .B(n3758), .ZN(n3760) );
  NAND2_X1 U4529 ( .A1(n3760), .A2(n3883), .ZN(n3764) );
  NOR2_X1 U4530 ( .A1(STATE_REG_SCAN_IN), .A2(n2790), .ZN(n4627) );
  AOI21_X1 U4531 ( .B1(n3885), .B2(n4370), .A(n4627), .ZN(n3763) );
  AOI22_X1 U4532 ( .A1(n4383), .A2(n3887), .B1(n3886), .B2(n4057), .ZN(n3762)
         );
  NAND2_X1 U4533 ( .A1(n3890), .A2(n4377), .ZN(n3761) );
  NAND4_X1 U4534 ( .A1(n3764), .A2(n3763), .A3(n3762), .A4(n3761), .ZN(U3225)
         );
  INV_X1 U4535 ( .A(n3765), .ZN(n3766) );
  NOR2_X1 U4536 ( .A1(n3767), .A2(n3766), .ZN(n3769) );
  XNOR2_X1 U4537 ( .A(n3769), .B(n3768), .ZN(n3770) );
  NAND2_X1 U4538 ( .A1(n3770), .A2(n3883), .ZN(n3775) );
  AOI22_X1 U4539 ( .A1(n3885), .A2(n4192), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3774) );
  AOI22_X1 U4540 ( .A1(n4237), .A2(n3887), .B1(n3886), .B2(n4054), .ZN(n3773)
         );
  INV_X1 U4541 ( .A(n3771), .ZN(n4234) );
  NAND2_X1 U4542 ( .A1(n3890), .A2(n4234), .ZN(n3772) );
  NAND4_X1 U4543 ( .A1(n3775), .A2(n3774), .A3(n3773), .A4(n3772), .ZN(U3226)
         );
  AOI21_X1 U4544 ( .B1(n3776), .B2(n3777), .A(n3829), .ZN(n3779) );
  NAND2_X1 U4545 ( .A1(n3779), .A2(n3778), .ZN(n3786) );
  AOI21_X1 U4546 ( .B1(n3885), .B2(n4068), .A(n3780), .ZN(n3785) );
  AOI22_X1 U4547 ( .A1(n3781), .A2(n3887), .B1(n3886), .B2(n2592), .ZN(n3784)
         );
  NAND2_X1 U4548 ( .A1(n3890), .A2(n3782), .ZN(n3783) );
  NAND4_X1 U4549 ( .A1(n3786), .A2(n3785), .A3(n3784), .A4(n3783), .ZN(U3227)
         );
  XNOR2_X1 U4550 ( .A(n3787), .B(n3788), .ZN(n3789) );
  NAND2_X1 U4551 ( .A1(n3789), .A2(n3883), .ZN(n3795) );
  INV_X1 U4552 ( .A(REG3_REG_9__SCAN_IN), .ZN(n4870) );
  NOR2_X1 U4553 ( .A1(STATE_REG_SCAN_IN), .A2(n4870), .ZN(n4564) );
  AOI21_X1 U4554 ( .B1(n3885), .B2(n4063), .A(n4564), .ZN(n3794) );
  AOI22_X1 U4555 ( .A1(n3790), .A2(n3887), .B1(n3886), .B2(n4065), .ZN(n3793)
         );
  NAND2_X1 U4556 ( .A1(n3890), .A2(n3791), .ZN(n3792) );
  NAND4_X1 U4557 ( .A1(n3795), .A2(n3794), .A3(n3793), .A4(n3792), .ZN(U3228)
         );
  INV_X1 U4558 ( .A(n3796), .ZN(n3798) );
  NAND2_X1 U4559 ( .A1(n3798), .A2(n3797), .ZN(n3799) );
  XNOR2_X1 U4560 ( .A(n3800), .B(n3799), .ZN(n3801) );
  NAND2_X1 U4561 ( .A1(n3801), .A2(n3883), .ZN(n3806) );
  AOI22_X1 U4562 ( .A1(n3885), .A2(n4273), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3805) );
  AOI22_X1 U4563 ( .A1(n4306), .A2(n3887), .B1(n3886), .B2(n4350), .ZN(n3804)
         );
  NAND2_X1 U4564 ( .A1(n3890), .A2(n3802), .ZN(n3803) );
  NAND4_X1 U4565 ( .A1(n3806), .A2(n3805), .A3(n3804), .A4(n3803), .ZN(U3230)
         );
  XNOR2_X1 U4566 ( .A(n3808), .B(n3807), .ZN(n3809) );
  XNOR2_X1 U4567 ( .A(n3810), .B(n3809), .ZN(n3811) );
  NAND2_X1 U4568 ( .A1(n3811), .A2(n3883), .ZN(n3818) );
  AOI21_X1 U4569 ( .B1(n3886), .B2(n4061), .A(n3812), .ZN(n3817) );
  AOI22_X1 U4570 ( .A1(n3813), .A2(n3887), .B1(n3885), .B2(n4059), .ZN(n3816)
         );
  NAND2_X1 U4571 ( .A1(n3890), .A2(n3814), .ZN(n3815) );
  NAND4_X1 U4572 ( .A1(n3818), .A2(n3817), .A3(n3816), .A4(n3815), .ZN(U3231)
         );
  AOI21_X1 U4573 ( .B1(n3821), .B2(n3820), .A(n3819), .ZN(n3830) );
  OAI22_X1 U4574 ( .A1(n3823), .A2(n4425), .B1(STATE_REG_SCAN_IN), .B2(n3822), 
        .ZN(n3827) );
  OAI22_X1 U4575 ( .A1(n3825), .A2(n4276), .B1(n3824), .B2(n4308), .ZN(n3826)
         );
  AOI211_X1 U4576 ( .C1(n4277), .C2(n3890), .A(n3827), .B(n3826), .ZN(n3828)
         );
  OAI21_X1 U4577 ( .B1(n3830), .B2(n3829), .A(n3828), .ZN(U3232) );
  XNOR2_X1 U4578 ( .A(n3832), .B(n3831), .ZN(n3833) );
  XNOR2_X1 U4579 ( .A(n3834), .B(n3833), .ZN(n3835) );
  NAND2_X1 U4580 ( .A1(n3835), .A2(n3883), .ZN(n3842) );
  NOR2_X1 U4581 ( .A1(STATE_REG_SCAN_IN), .A2(n3836), .ZN(n4584) );
  AOI21_X1 U4582 ( .B1(n3885), .B2(n4061), .A(n4584), .ZN(n3841) );
  AOI22_X1 U4583 ( .A1(n3837), .A2(n3887), .B1(n3886), .B2(n4063), .ZN(n3840)
         );
  NAND2_X1 U4584 ( .A1(n3890), .A2(n3838), .ZN(n3839) );
  NAND4_X1 U4585 ( .A1(n3842), .A2(n3841), .A3(n3840), .A4(n3839), .ZN(U3233)
         );
  INV_X1 U4586 ( .A(n3846), .ZN(n3843) );
  NOR2_X1 U4587 ( .A1(n3844), .A2(n3843), .ZN(n3849) );
  AOI21_X1 U4588 ( .B1(n3847), .B2(n3846), .A(n3845), .ZN(n3848) );
  OAI21_X1 U4589 ( .B1(n3849), .B2(n3848), .A(n3883), .ZN(n3854) );
  NOR2_X1 U4590 ( .A1(n3850), .A2(STATE_REG_SCAN_IN), .ZN(n4111) );
  AOI21_X1 U4591 ( .B1(n3885), .B2(n4350), .A(n4111), .ZN(n3853) );
  AOI22_X1 U4592 ( .A1(n4349), .A2(n3887), .B1(n3886), .B2(n4056), .ZN(n3852)
         );
  NAND2_X1 U4593 ( .A1(n3890), .A2(n4358), .ZN(n3851) );
  NAND4_X1 U4594 ( .A1(n3854), .A2(n3853), .A3(n3852), .A4(n3851), .ZN(U3235)
         );
  XNOR2_X1 U4595 ( .A(n3856), .B(n3855), .ZN(n3857) );
  XNOR2_X1 U4596 ( .A(n3858), .B(n3857), .ZN(n3859) );
  NAND2_X1 U4597 ( .A1(n3859), .A2(n3883), .ZN(n3866) );
  AOI21_X1 U4598 ( .B1(n3885), .B2(n4066), .A(n3860), .ZN(n3865) );
  AOI22_X1 U4599 ( .A1(n3861), .A2(n3887), .B1(n3886), .B2(n4068), .ZN(n3864)
         );
  NAND2_X1 U4600 ( .A1(n3890), .A2(n3862), .ZN(n3863) );
  NAND4_X1 U4601 ( .A1(n3866), .A2(n3865), .A3(n3864), .A4(n3863), .ZN(U3236)
         );
  NOR2_X1 U4602 ( .A1(n2422), .A2(n3868), .ZN(n3869) );
  XNOR2_X1 U4603 ( .A(n3870), .B(n3869), .ZN(n3871) );
  NAND2_X1 U4604 ( .A1(n3871), .A2(n3883), .ZN(n3877) );
  AOI22_X1 U4605 ( .A1(n4400), .A2(n3885), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3876) );
  AOI22_X1 U4606 ( .A1(n3872), .A2(n3887), .B1(n3886), .B2(n4192), .ZN(n3875)
         );
  INV_X1 U4607 ( .A(n4200), .ZN(n3873) );
  NAND2_X1 U4608 ( .A1(n3890), .A2(n3873), .ZN(n3874) );
  NAND4_X1 U4609 ( .A1(n3877), .A2(n3876), .A3(n3875), .A4(n3874), .ZN(U3237)
         );
  INV_X1 U4610 ( .A(n3878), .ZN(n3880) );
  NAND2_X1 U4611 ( .A1(n3880), .A2(n3879), .ZN(n3882) );
  XNOR2_X1 U4612 ( .A(n3882), .B(n3881), .ZN(n3884) );
  NAND2_X1 U4613 ( .A1(n3884), .A2(n3883), .ZN(n3894) );
  AND2_X1 U4614 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4608) );
  AOI21_X1 U4615 ( .B1(n3885), .B2(n4057), .A(n4608), .ZN(n3893) );
  AOI22_X1 U4616 ( .A1(n3888), .A2(n3887), .B1(n3886), .B2(n4059), .ZN(n3892)
         );
  NAND2_X1 U4617 ( .A1(n3890), .A2(n3889), .ZN(n3891) );
  NAND4_X1 U4618 ( .A1(n3894), .A2(n3893), .A3(n3892), .A4(n3891), .ZN(U3238)
         );
  INV_X1 U4619 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4390) );
  NAND2_X1 U4620 ( .A1(n2840), .A2(REG2_REG_31__SCAN_IN), .ZN(n3897) );
  NAND2_X1 U4621 ( .A1(n3895), .A2(REG0_REG_31__SCAN_IN), .ZN(n3896) );
  OAI211_X1 U4622 ( .C1(n2564), .C2(n4390), .A(n3897), .B(n3896), .ZN(n4151)
         );
  NAND2_X1 U4623 ( .A1(n2552), .A2(DATAI_31_), .ZN(n4152) );
  NAND2_X1 U4624 ( .A1(n2552), .A2(DATAI_30_), .ZN(n4148) );
  NAND2_X1 U4625 ( .A1(n4053), .A2(n4148), .ZN(n4037) );
  OAI21_X1 U4626 ( .B1(n4151), .B2(n4152), .A(n4037), .ZN(n4006) );
  INV_X1 U4627 ( .A(n4006), .ZN(n4044) );
  XNOR2_X1 U4628 ( .A(n4054), .B(n4260), .ZN(n4242) );
  INV_X1 U4629 ( .A(n4242), .ZN(n4252) );
  NAND2_X1 U4630 ( .A1(n2358), .A2(n4671), .ZN(n3898) );
  NOR4_X1 U4631 ( .A1(n4177), .A2(n3899), .A3(n4252), .A4(n3898), .ZN(n3909)
         );
  OR2_X1 U4632 ( .A1(n4186), .A2(n2301), .ZN(n4207) );
  INV_X1 U4633 ( .A(n4207), .ZN(n4208) );
  INV_X1 U4634 ( .A(n3986), .ZN(n3901) );
  NAND4_X1 U4635 ( .A1(n4285), .A2(n3904), .A3(n3903), .A4(n3902), .ZN(n3907)
         );
  NOR4_X1 U4636 ( .A1(n4195), .A2(n3907), .A3(n3906), .A4(n3905), .ZN(n3908)
         );
  NAND4_X1 U4637 ( .A1(n3909), .A2(n4161), .A3(n4208), .A4(n3908), .ZN(n3929)
         );
  XNOR2_X1 U4638 ( .A(n4350), .B(n4336), .ZN(n4330) );
  NOR4_X1 U4639 ( .A1(n3057), .A2(n3911), .A3(n3056), .A4(n3910), .ZN(n3926)
         );
  NAND2_X1 U4640 ( .A1(n2256), .A2(n3912), .ZN(n4229) );
  INV_X1 U4641 ( .A(n3913), .ZN(n3915) );
  OR2_X1 U4642 ( .A1(n3915), .A2(n3914), .ZN(n4304) );
  INV_X1 U4643 ( .A(n4304), .ZN(n3916) );
  NAND2_X1 U4644 ( .A1(n4151), .A2(n4152), .ZN(n4007) );
  OAI21_X1 U4645 ( .B1(n4053), .B2(n4148), .A(n4007), .ZN(n3999) );
  NOR4_X1 U4646 ( .A1(n4229), .A2(n3916), .A3(n4539), .A4(n3999), .ZN(n3925)
         );
  NAND2_X1 U4647 ( .A1(n4324), .A2(n4244), .ZN(n4365) );
  NOR4_X1 U4648 ( .A1(n4365), .A2(n3919), .A3(n3918), .A4(n3917), .ZN(n3924)
         );
  NOR4_X1 U4649 ( .A1(n4348), .A2(n3922), .A3(n3921), .A4(n3920), .ZN(n3923)
         );
  NAND4_X1 U4650 ( .A1(n3926), .A2(n3925), .A3(n3924), .A4(n3923), .ZN(n3927)
         );
  NOR4_X1 U4651 ( .A1(n3929), .A2(n4330), .A3(n3928), .A4(n3927), .ZN(n3998)
         );
  AND2_X1 U4652 ( .A1(n2256), .A2(n3930), .ZN(n4008) );
  INV_X1 U4653 ( .A(n3931), .ZN(n3934) );
  OAI211_X1 U4654 ( .C1(n3934), .C2(n4539), .A(n3933), .B(n3932), .ZN(n3937)
         );
  NAND3_X1 U4655 ( .A1(n3937), .A2(n3936), .A3(n3935), .ZN(n3940) );
  NAND3_X1 U4656 ( .A1(n3940), .A2(n3939), .A3(n3938), .ZN(n3943) );
  NAND3_X1 U4657 ( .A1(n3943), .A2(n3942), .A3(n3941), .ZN(n3946) );
  NAND4_X1 U4658 ( .A1(n3946), .A2(n3945), .A3(n3944), .A4(n3959), .ZN(n3949)
         );
  NAND3_X1 U4659 ( .A1(n3949), .A2(n3948), .A3(n3947), .ZN(n3956) );
  AND2_X1 U4660 ( .A1(n3951), .A2(n3950), .ZN(n3960) );
  INV_X1 U4661 ( .A(n3952), .ZN(n3955) );
  INV_X1 U4662 ( .A(n3953), .ZN(n3954) );
  AOI211_X1 U4663 ( .C1(n3956), .C2(n3960), .A(n3955), .B(n3954), .ZN(n3968)
         );
  NAND2_X1 U4664 ( .A1(n3958), .A2(n3957), .ZN(n3967) );
  INV_X1 U4665 ( .A(n3959), .ZN(n3963) );
  INV_X1 U4666 ( .A(n3960), .ZN(n3962) );
  NOR3_X1 U4667 ( .A1(n3963), .A2(n3962), .A3(n3961), .ZN(n3965) );
  INV_X1 U4668 ( .A(n3970), .ZN(n3964) );
  NAND2_X1 U4669 ( .A1(n3967), .A2(n3976), .ZN(n4009) );
  OAI21_X1 U4670 ( .B1(n3965), .B2(n3964), .A(n4009), .ZN(n3966) );
  OAI21_X1 U4671 ( .B1(n3968), .B2(n3967), .A(n3966), .ZN(n3974) );
  NAND2_X1 U4672 ( .A1(n3970), .A2(n3969), .ZN(n3971) );
  NAND4_X1 U4673 ( .A1(n3974), .A2(n3973), .A3(n3972), .A4(n3971), .ZN(n3981)
         );
  INV_X1 U4674 ( .A(n3975), .ZN(n3978) );
  NAND2_X1 U4675 ( .A1(n3977), .A2(n3976), .ZN(n4010) );
  OAI21_X1 U4676 ( .B1(n3978), .B2(n4010), .A(n4009), .ZN(n3980) );
  INV_X1 U4677 ( .A(n3979), .ZN(n4012) );
  AOI21_X1 U4678 ( .B1(n3981), .B2(n3980), .A(n4012), .ZN(n3985) );
  INV_X1 U4679 ( .A(n4013), .ZN(n3984) );
  INV_X1 U4680 ( .A(n3982), .ZN(n3983) );
  OAI21_X1 U4681 ( .B1(n3985), .B2(n3984), .A(n3983), .ZN(n3987) );
  AOI211_X1 U4682 ( .C1(n3987), .C2(n4249), .A(n3986), .B(n4248), .ZN(n3988)
         );
  NOR2_X1 U4683 ( .A1(n3988), .A2(n4020), .ZN(n3990) );
  OAI21_X1 U4684 ( .B1(n3990), .B2(n3989), .A(n4024), .ZN(n3991) );
  NAND2_X1 U4685 ( .A1(n4008), .A2(n3991), .ZN(n3996) );
  INV_X1 U4686 ( .A(n4163), .ZN(n4001) );
  OAI21_X1 U4687 ( .B1(n4000), .B2(n4001), .A(n3992), .ZN(n4002) );
  NOR2_X1 U4688 ( .A1(n3993), .A2(n4002), .ZN(n4032) );
  INV_X1 U4689 ( .A(n4032), .ZN(n3994) );
  AOI211_X1 U4690 ( .C1(n4022), .C2(n3996), .A(n3995), .B(n3994), .ZN(n3997)
         );
  MUX2_X1 U4691 ( .A(n3998), .B(n3997), .S(n2506), .Z(n4043) );
  NOR2_X1 U4692 ( .A1(n4029), .A2(n4028), .ZN(n4003) );
  AOI21_X1 U4693 ( .B1(n4001), .B2(n4000), .A(n3999), .ZN(n4026) );
  OAI21_X1 U4694 ( .B1(n4003), .B2(n4002), .A(n4026), .ZN(n4031) );
  INV_X1 U4695 ( .A(n4031), .ZN(n4004) );
  AOI211_X1 U4696 ( .C1(n4007), .C2(n4006), .A(n4005), .B(n4004), .ZN(n4042)
         );
  INV_X1 U4697 ( .A(n4008), .ZN(n4025) );
  OAI21_X1 U4698 ( .B1(n4011), .B2(n4010), .A(n4009), .ZN(n4014) );
  AOI21_X1 U4699 ( .B1(n4014), .B2(n4013), .A(n4012), .ZN(n4017) );
  INV_X1 U4700 ( .A(n4249), .ZN(n4016) );
  OAI21_X1 U4701 ( .B1(n4017), .B2(n4016), .A(n4015), .ZN(n4018) );
  INV_X1 U4702 ( .A(n4018), .ZN(n4021) );
  OAI21_X1 U4703 ( .B1(n4021), .B2(n4020), .A(n4019), .ZN(n4023) );
  OAI221_X1 U4704 ( .B1(n4025), .B2(n4024), .C1(n4025), .C2(n4023), .A(n4022), 
        .ZN(n4030) );
  INV_X1 U4705 ( .A(n4026), .ZN(n4027) );
  NOR4_X1 U4706 ( .A1(n4030), .A2(n4029), .A3(n4028), .A4(n4027), .ZN(n4035)
         );
  INV_X1 U4707 ( .A(n4177), .ZN(n4033) );
  AOI21_X1 U4708 ( .B1(n4033), .B2(n4032), .A(n4031), .ZN(n4034) );
  OAI22_X1 U4709 ( .A1(n4035), .A2(n4034), .B1(n4151), .B2(n4148), .ZN(n4036)
         );
  INV_X1 U4710 ( .A(n4036), .ZN(n4040) );
  AOI21_X1 U4711 ( .B1(n4037), .B2(n4151), .A(n4152), .ZN(n4039) );
  NOR3_X1 U4712 ( .A1(n4040), .A2(n4039), .A3(n4038), .ZN(n4041) );
  AOI211_X1 U4713 ( .C1(n4044), .C2(n4043), .A(n4042), .B(n4041), .ZN(n4045)
         );
  XNOR2_X1 U4714 ( .A(n4045), .B(n4144), .ZN(n4052) );
  NOR2_X1 U4715 ( .A1(n4047), .A2(n4046), .ZN(n4050) );
  OAI21_X1 U4716 ( .B1(n4051), .B2(n4048), .A(B_REG_SCAN_IN), .ZN(n4049) );
  OAI22_X1 U4717 ( .A1(n4052), .A2(n4051), .B1(n4050), .B2(n4049), .ZN(U3239)
         );
  MUX2_X1 U4718 ( .A(n4151), .B(DATAO_REG_31__SCAN_IN), .S(n4071), .Z(U3581)
         );
  MUX2_X1 U4719 ( .A(n4053), .B(DATAO_REG_30__SCAN_IN), .S(n4071), .Z(U3580)
         );
  MUX2_X1 U4720 ( .A(n4163), .B(DATAO_REG_29__SCAN_IN), .S(n4071), .Z(U3579)
         );
  MUX2_X1 U4721 ( .A(n4179), .B(DATAO_REG_28__SCAN_IN), .S(n4071), .Z(U3578)
         );
  MUX2_X1 U4722 ( .A(DATAO_REG_27__SCAN_IN), .B(n4400), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4723 ( .A(n4409), .B(DATAO_REG_26__SCAN_IN), .S(n4071), .Z(U3576)
         );
  MUX2_X1 U4724 ( .A(DATAO_REG_25__SCAN_IN), .B(n4192), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4725 ( .A(n4212), .B(DATAO_REG_24__SCAN_IN), .S(n4071), .Z(U3574)
         );
  MUX2_X1 U4726 ( .A(n4054), .B(DATAO_REG_23__SCAN_IN), .S(n4071), .Z(U3573)
         );
  MUX2_X1 U4727 ( .A(DATAO_REG_22__SCAN_IN), .B(n4257), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4728 ( .A(n4273), .B(DATAO_REG_21__SCAN_IN), .S(n4071), .Z(U3571)
         );
  MUX2_X1 U4729 ( .A(n4055), .B(DATAO_REG_20__SCAN_IN), .S(n4071), .Z(U3570)
         );
  MUX2_X1 U4730 ( .A(n4350), .B(DATAO_REG_19__SCAN_IN), .S(n4071), .Z(U3569)
         );
  MUX2_X1 U4731 ( .A(n4370), .B(DATAO_REG_18__SCAN_IN), .S(n4071), .Z(U3568)
         );
  MUX2_X1 U4732 ( .A(n4056), .B(DATAO_REG_17__SCAN_IN), .S(n4071), .Z(U3567)
         );
  MUX2_X1 U4733 ( .A(n4057), .B(DATAO_REG_16__SCAN_IN), .S(n4071), .Z(U3566)
         );
  MUX2_X1 U4734 ( .A(n4058), .B(DATAO_REG_15__SCAN_IN), .S(n4071), .Z(U3565)
         );
  MUX2_X1 U4735 ( .A(n4059), .B(DATAO_REG_14__SCAN_IN), .S(n4071), .Z(U3564)
         );
  MUX2_X1 U4736 ( .A(n4060), .B(DATAO_REG_13__SCAN_IN), .S(n4071), .Z(U3563)
         );
  MUX2_X1 U4737 ( .A(n4061), .B(DATAO_REG_12__SCAN_IN), .S(n4071), .Z(U3562)
         );
  MUX2_X1 U4738 ( .A(n4062), .B(DATAO_REG_11__SCAN_IN), .S(n4071), .Z(U3561)
         );
  MUX2_X1 U4739 ( .A(n4063), .B(DATAO_REG_10__SCAN_IN), .S(n4071), .Z(U3560)
         );
  MUX2_X1 U4740 ( .A(n4064), .B(DATAO_REG_9__SCAN_IN), .S(n4071), .Z(U3559) );
  MUX2_X1 U4741 ( .A(n4065), .B(DATAO_REG_8__SCAN_IN), .S(n4071), .Z(U3558) );
  MUX2_X1 U4742 ( .A(n4066), .B(DATAO_REG_7__SCAN_IN), .S(n4071), .Z(U3557) );
  MUX2_X1 U4743 ( .A(n4067), .B(DATAO_REG_6__SCAN_IN), .S(n4071), .Z(U3556) );
  MUX2_X1 U4744 ( .A(n4068), .B(DATAO_REG_5__SCAN_IN), .S(n4071), .Z(U3555) );
  MUX2_X1 U4745 ( .A(n4069), .B(DATAO_REG_4__SCAN_IN), .S(n4071), .Z(U3554) );
  MUX2_X1 U4746 ( .A(n2592), .B(DATAO_REG_3__SCAN_IN), .S(n4071), .Z(U3553) );
  MUX2_X1 U4747 ( .A(n2574), .B(DATAO_REG_2__SCAN_IN), .S(n4071), .Z(U3552) );
  MUX2_X1 U4748 ( .A(n4070), .B(DATAO_REG_1__SCAN_IN), .S(n4071), .Z(U3551) );
  MUX2_X1 U4749 ( .A(n4072), .B(DATAO_REG_0__SCAN_IN), .S(n4071), .Z(U3550) );
  INV_X1 U4750 ( .A(n4073), .ZN(n4075) );
  AOI21_X1 U4751 ( .B1(n2530), .B2(n4074), .A(n4075), .ZN(n4076) );
  MUX2_X1 U4752 ( .A(n4076), .B(n4075), .S(IR_REG_0__SCAN_IN), .Z(n4078) );
  AOI22_X1 U4753 ( .A1(n4078), .A2(n4077), .B1(REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4081) );
  NAND3_X1 U4754 ( .A1(n4629), .A2(IR_REG_0__SCAN_IN), .A3(n2530), .ZN(n4080)
         );
  NAND2_X1 U4755 ( .A1(n4628), .A2(ADDR_REG_0__SCAN_IN), .ZN(n4079) );
  NAND3_X1 U4756 ( .A1(n4081), .A2(n4080), .A3(n4079), .ZN(U3240) );
  NAND2_X1 U4757 ( .A1(n4092), .A2(n4549), .ZN(n4091) );
  OAI211_X1 U4758 ( .C1(n2236), .C2(n4084), .A(n4587), .B(n4083), .ZN(n4090)
         );
  OAI211_X1 U4759 ( .C1(n4087), .C2(n4086), .A(n4629), .B(n4085), .ZN(n4089)
         );
  AOI22_X1 U4760 ( .A1(n4628), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4088) );
  NAND4_X1 U4761 ( .A1(n4091), .A2(n4090), .A3(n4089), .A4(n4088), .ZN(U3241)
         );
  NAND2_X1 U4762 ( .A1(n4092), .A2(n4547), .ZN(n4101) );
  OAI211_X1 U4763 ( .C1(REG1_REG_3__SCAN_IN), .C2(n4094), .A(n4629), .B(n4093), 
        .ZN(n4100) );
  AOI22_X1 U4764 ( .A1(n4628), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n4099) );
  XNOR2_X1 U4765 ( .A(n4096), .B(n4095), .ZN(n4097) );
  NAND2_X1 U4766 ( .A1(n4587), .A2(n4097), .ZN(n4098) );
  NAND4_X1 U4767 ( .A1(n4101), .A2(n4100), .A3(n4099), .A4(n4098), .ZN(U3243)
         );
  XOR2_X1 U4768 ( .A(REG1_REG_18__SCAN_IN), .B(n4138), .Z(n4139) );
  NOR2_X1 U4769 ( .A1(n4127), .A2(REG1_REG_17__SCAN_IN), .ZN(n4110) );
  NAND2_X1 U4770 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4123), .ZN(n4107) );
  INV_X1 U4771 ( .A(n4123), .ZN(n4664) );
  AOI22_X1 U4772 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4123), .B1(n4664), .B2(
        n3602), .ZN(n4611) );
  INV_X1 U4773 ( .A(n4102), .ZN(n4104) );
  NAND2_X1 U4774 ( .A1(n4104), .A2(n4103), .ZN(n4105) );
  NAND2_X1 U4775 ( .A1(n4120), .A2(n4105), .ZN(n4106) );
  XNOR2_X1 U4776 ( .A(n4105), .B(n2336), .ZN(n4602) );
  NAND2_X1 U4777 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4602), .ZN(n4601) );
  NAND2_X1 U4778 ( .A1(n4106), .A2(n4601), .ZN(n4610) );
  NAND2_X1 U4779 ( .A1(n4611), .A2(n4610), .ZN(n4609) );
  NOR2_X1 U4780 ( .A1(n4124), .A2(n4108), .ZN(n4109) );
  INV_X1 U4781 ( .A(n4124), .ZN(n4663) );
  AOI22_X1 U4782 ( .A1(n4127), .A2(n4465), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4662), .ZN(n4630) );
  NOR2_X1 U4783 ( .A1(n4631), .A2(n4630), .ZN(n4632) );
  XOR2_X1 U4784 ( .A(n4139), .B(n4140), .Z(n4132) );
  INV_X1 U4785 ( .A(n4138), .ZN(n4113) );
  AOI21_X1 U4786 ( .B1(n4628), .B2(ADDR_REG_18__SCAN_IN), .A(n4111), .ZN(n4112) );
  OAI21_X1 U4787 ( .B1(n4635), .B2(n4113), .A(n4112), .ZN(n4131) );
  INV_X1 U4788 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4115) );
  NOR2_X1 U4789 ( .A1(n4138), .A2(n4115), .ZN(n4114) );
  AOI21_X1 U4790 ( .B1(n4138), .B2(n4115), .A(n4114), .ZN(n4129) );
  NOR2_X1 U4791 ( .A1(n4127), .A2(REG2_REG_17__SCAN_IN), .ZN(n4116) );
  AOI21_X1 U4792 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4127), .A(n4116), .ZN(n4625) );
  NOR2_X1 U4793 ( .A1(n2336), .A2(n4119), .ZN(n4121) );
  INV_X1 U4794 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4598) );
  NAND2_X1 U4795 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4123), .ZN(n4122) );
  OAI21_X1 U4796 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4123), .A(n4122), .ZN(n4605) );
  NAND2_X1 U4797 ( .A1(n4125), .A2(n4663), .ZN(n4126) );
  XNOR2_X1 U4798 ( .A(n4125), .B(n4124), .ZN(n4615) );
  NAND2_X1 U4799 ( .A1(n4615), .A2(n3610), .ZN(n4614) );
  NAND2_X1 U4800 ( .A1(n4126), .A2(n4614), .ZN(n4623) );
  NAND2_X1 U4801 ( .A1(n4625), .A2(n4623), .ZN(n4624) );
  AOI211_X1 U4802 ( .C1(n4129), .C2(n4128), .A(n4135), .B(n4622), .ZN(n4130)
         );
  AOI211_X1 U4803 ( .C1(n4132), .C2(n4629), .A(n4131), .B(n4130), .ZN(n4133)
         );
  INV_X1 U4804 ( .A(n4133), .ZN(U3258) );
  INV_X1 U4805 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4134) );
  MUX2_X1 U4806 ( .A(REG2_REG_19__SCAN_IN), .B(n4134), .S(n4540), .Z(n4136) );
  INV_X1 U4807 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4137) );
  MUX2_X1 U4808 ( .A(n4137), .B(REG1_REG_19__SCAN_IN), .S(n4540), .Z(n4141) );
  NAND2_X1 U4809 ( .A1(n4628), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4142) );
  OAI211_X1 U4810 ( .C1(n4635), .C2(n4144), .A(n4143), .B(n4142), .ZN(n4145)
         );
  OAI21_X1 U4811 ( .B1(n4147), .B2(n4622), .A(n4146), .ZN(U3259) );
  XNOR2_X1 U4812 ( .A(n4393), .B(n4152), .ZN(n4483) );
  INV_X1 U4813 ( .A(n4149), .ZN(n4150) );
  NAND2_X1 U4814 ( .A1(n4151), .A2(n4150), .ZN(n4397) );
  OAI21_X1 U4815 ( .B1(n4152), .B2(n4459), .A(n4397), .ZN(n4480) );
  NAND2_X1 U4816 ( .A1(n4648), .A2(n4480), .ZN(n4154) );
  NAND2_X1 U4817 ( .A1(n4378), .A2(REG2_REG_31__SCAN_IN), .ZN(n4153) );
  OAI211_X1 U4818 ( .C1(n4483), .C2(n4385), .A(n4154), .B(n4153), .ZN(U3260)
         );
  XNOR2_X1 U4819 ( .A(n4155), .B(n4161), .ZN(n4403) );
  OAI21_X1 U4820 ( .B1(n4172), .B2(n4157), .A(n4156), .ZN(n4490) );
  INV_X1 U4821 ( .A(n4490), .ZN(n4167) );
  AOI22_X1 U4822 ( .A1(n4158), .A2(n4636), .B1(n4378), .B2(
        REG2_REG_28__SCAN_IN), .ZN(n4160) );
  NAND2_X1 U4823 ( .A1(n4382), .A2(n2324), .ZN(n4159) );
  OAI211_X1 U4824 ( .C1(n4185), .C2(n4380), .A(n4160), .B(n4159), .ZN(n4166)
         );
  XNOR2_X1 U4825 ( .A(n4162), .B(n4161), .ZN(n4164) );
  AOI22_X1 U4826 ( .A1(n4164), .A2(n4367), .B1(n4369), .B2(n4163), .ZN(n4402)
         );
  NOR2_X1 U4827 ( .A1(n4402), .A2(n4378), .ZN(n4165) );
  AOI211_X1 U4828 ( .C1(n4652), .C2(n4167), .A(n4166), .B(n4165), .ZN(n4168)
         );
  OAI21_X1 U4829 ( .B1(n4403), .B2(n4388), .A(n4168), .ZN(U3262) );
  XNOR2_X1 U4830 ( .A(n4169), .B(n4177), .ZN(n4412) );
  NOR2_X1 U4831 ( .A1(n4197), .A2(n4170), .ZN(n4171) );
  INV_X1 U4832 ( .A(n4494), .ZN(n4183) );
  INV_X1 U4833 ( .A(n4409), .ZN(n4176) );
  AOI22_X1 U4834 ( .A1(n4378), .A2(REG2_REG_27__SCAN_IN), .B1(n4173), .B2(
        n4636), .ZN(n4175) );
  NAND2_X1 U4835 ( .A1(n4382), .A2(n4407), .ZN(n4174) );
  OAI211_X1 U4836 ( .C1(n4176), .C2(n4380), .A(n4175), .B(n4174), .ZN(n4182)
         );
  XNOR2_X1 U4837 ( .A(n4178), .B(n4177), .ZN(n4180) );
  AOI22_X1 U4838 ( .A1(n4180), .A2(n4367), .B1(n4369), .B2(n4179), .ZN(n4411)
         );
  NOR2_X1 U4839 ( .A1(n4411), .A2(n4378), .ZN(n4181) );
  AOI211_X1 U4840 ( .C1(n4652), .C2(n4183), .A(n4182), .B(n4181), .ZN(n4184)
         );
  OAI21_X1 U4841 ( .B1(n4412), .B2(n4388), .A(n4184), .ZN(U3263) );
  OAI22_X1 U4842 ( .A1(n4185), .A2(n4331), .B1(n4459), .B2(n4199), .ZN(n4191)
         );
  NOR2_X1 U4843 ( .A1(n4187), .A2(n4186), .ZN(n4188) );
  XOR2_X1 U4844 ( .A(n4195), .B(n4188), .Z(n4189) );
  NOR2_X1 U4845 ( .A1(n4189), .A2(n4334), .ZN(n4190) );
  AOI211_X1 U4846 ( .C1(n4408), .C2(n4192), .A(n4191), .B(n4190), .ZN(n4415)
         );
  XOR2_X1 U4848 ( .A(n4195), .B(n4194), .Z(n4417) );
  NAND2_X1 U4849 ( .A1(n4417), .A2(n4196), .ZN(n4205) );
  INV_X1 U4850 ( .A(n4197), .ZN(n4198) );
  OAI21_X1 U4851 ( .B1(n4217), .B2(n4199), .A(n4198), .ZN(n4498) );
  INV_X1 U4852 ( .A(n4498), .ZN(n4203) );
  INV_X1 U4853 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4201) );
  OAI22_X1 U4854 ( .A1(n4648), .A2(n4201), .B1(n4200), .B2(n4645), .ZN(n4202)
         );
  AOI21_X1 U4855 ( .B1(n4203), .B2(n4652), .A(n4202), .ZN(n4204) );
  OAI211_X1 U4856 ( .C1(n4378), .C2(n4415), .A(n4205), .B(n4204), .ZN(U3264)
         );
  XOR2_X1 U4857 ( .A(n4207), .B(n4206), .Z(n4421) );
  INV_X1 U4858 ( .A(n4421), .ZN(n4225) );
  XNOR2_X1 U4859 ( .A(n4209), .B(n4208), .ZN(n4210) );
  NAND2_X1 U4860 ( .A1(n4210), .A2(n4367), .ZN(n4216) );
  NAND2_X1 U4861 ( .A1(n4409), .A2(n4369), .ZN(n4214) );
  AOI22_X1 U4862 ( .A1(n4212), .A2(n4408), .B1(n4211), .B2(n4406), .ZN(n4213)
         );
  AND2_X1 U4863 ( .A1(n4214), .A2(n4213), .ZN(n4215) );
  NAND2_X1 U4864 ( .A1(n4216), .A2(n4215), .ZN(n4420) );
  INV_X1 U4865 ( .A(n4233), .ZN(n4220) );
  INV_X1 U4866 ( .A(n4217), .ZN(n4218) );
  OAI21_X1 U4867 ( .B1(n4220), .B2(n4219), .A(n4218), .ZN(n4502) );
  AOI22_X1 U4868 ( .A1(n4378), .A2(REG2_REG_25__SCAN_IN), .B1(n4221), .B2(
        n4636), .ZN(n4222) );
  OAI21_X1 U4869 ( .B1(n4502), .B2(n4385), .A(n4222), .ZN(n4223) );
  AOI21_X1 U4870 ( .B1(n4420), .B2(n4648), .A(n4223), .ZN(n4224) );
  OAI21_X1 U4871 ( .B1(n4225), .B2(n4388), .A(n4224), .ZN(U3265) );
  XNOR2_X1 U4872 ( .A(n4226), .B(n4229), .ZN(n4428) );
  INV_X1 U4873 ( .A(n4428), .ZN(n4241) );
  NAND2_X1 U4874 ( .A1(n4228), .A2(n4227), .ZN(n4230) );
  XNOR2_X1 U4875 ( .A(n4230), .B(n4229), .ZN(n4232) );
  OAI22_X1 U4876 ( .A1(n4232), .A2(n4334), .B1(n4231), .B2(n4331), .ZN(n4427)
         );
  OAI21_X1 U4877 ( .B1(n2318), .B2(n4424), .A(n4233), .ZN(n4506) );
  AOI22_X1 U4878 ( .A1(n4378), .A2(REG2_REG_24__SCAN_IN), .B1(n4234), .B2(
        n4636), .ZN(n4235) );
  OAI21_X1 U4879 ( .B1(n4425), .B2(n4380), .A(n4235), .ZN(n4236) );
  AOI21_X1 U4880 ( .B1(n4237), .B2(n4382), .A(n4236), .ZN(n4238) );
  OAI21_X1 U4881 ( .B1(n4506), .B2(n4385), .A(n4238), .ZN(n4239) );
  AOI21_X1 U4882 ( .B1(n4427), .B2(n4648), .A(n4239), .ZN(n4240) );
  OAI21_X1 U4883 ( .B1(n4241), .B2(n4388), .A(n4240), .ZN(U3266) );
  XNOR2_X1 U4884 ( .A(n4243), .B(n4242), .ZN(n4432) );
  INV_X1 U4885 ( .A(n4432), .ZN(n4267) );
  INV_X1 U4886 ( .A(n4244), .ZN(n4245) );
  INV_X1 U4887 ( .A(n4246), .ZN(n4247) );
  AOI21_X1 U4888 ( .B1(n4303), .B2(n4249), .A(n4248), .ZN(n4286) );
  NAND2_X1 U4889 ( .A1(n4286), .A2(n4285), .ZN(n4284) );
  OAI21_X1 U4890 ( .B1(n4270), .B2(n4271), .A(n4251), .ZN(n4253) );
  XNOR2_X1 U4891 ( .A(n4253), .B(n4252), .ZN(n4259) );
  OAI22_X1 U4892 ( .A1(n4255), .A2(n4331), .B1(n4459), .B2(n4254), .ZN(n4256)
         );
  AOI21_X1 U4893 ( .B1(n4408), .B2(n4257), .A(n4256), .ZN(n4258) );
  OAI21_X1 U4894 ( .B1(n4259), .B2(n4334), .A(n4258), .ZN(n4431) );
  NAND2_X1 U4895 ( .A1(n2244), .A2(n4260), .ZN(n4261) );
  NAND2_X1 U4896 ( .A1(n4262), .A2(n4261), .ZN(n4510) );
  AOI22_X1 U4897 ( .A1(n4378), .A2(REG2_REG_23__SCAN_IN), .B1(n4263), .B2(
        n4636), .ZN(n4264) );
  OAI21_X1 U4898 ( .B1(n4510), .B2(n4385), .A(n4264), .ZN(n4265) );
  AOI21_X1 U4899 ( .B1(n4431), .B2(n4648), .A(n4265), .ZN(n4266) );
  OAI21_X1 U4900 ( .B1(n4267), .B2(n4388), .A(n4266), .ZN(U3267) );
  OAI21_X1 U4901 ( .B1(n4269), .B2(n4271), .A(n4268), .ZN(n4435) );
  XOR2_X1 U4902 ( .A(n4271), .B(n4270), .Z(n4275) );
  OAI22_X1 U4903 ( .A1(n4425), .A2(n4331), .B1(n4276), .B2(n4459), .ZN(n4272)
         );
  AOI21_X1 U4904 ( .B1(n4408), .B2(n4273), .A(n4272), .ZN(n4274) );
  OAI21_X1 U4905 ( .B1(n4275), .B2(n4334), .A(n4274), .ZN(n4436) );
  OAI21_X1 U4906 ( .B1(n4291), .B2(n4276), .A(n2244), .ZN(n4514) );
  NOR2_X1 U4907 ( .A1(n4514), .A2(n4385), .ZN(n4281) );
  INV_X1 U4908 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4279) );
  INV_X1 U4909 ( .A(n4277), .ZN(n4278) );
  OAI22_X1 U4910 ( .A1(n4648), .A2(n4279), .B1(n4278), .B2(n4645), .ZN(n4280)
         );
  AOI211_X1 U4911 ( .C1(n4436), .C2(n4648), .A(n4281), .B(n4280), .ZN(n4282)
         );
  OAI21_X1 U4912 ( .B1(n4435), .B2(n4388), .A(n4282), .ZN(U3268) );
  XNOR2_X1 U4913 ( .A(n4283), .B(n4285), .ZN(n4444) );
  INV_X1 U4914 ( .A(n4444), .ZN(n4300) );
  OAI21_X1 U4915 ( .B1(n4286), .B2(n4285), .A(n4284), .ZN(n4287) );
  NAND2_X1 U4916 ( .A1(n4287), .A2(n4367), .ZN(n4290) );
  OR2_X1 U4917 ( .A1(n4288), .A2(n4331), .ZN(n4289) );
  NAND2_X1 U4918 ( .A1(n4290), .A2(n4289), .ZN(n4443) );
  INV_X1 U4919 ( .A(n4291), .ZN(n4292) );
  OAI21_X1 U4920 ( .B1(n2317), .B2(n4440), .A(n4292), .ZN(n4518) );
  AOI22_X1 U4921 ( .A1(n4378), .A2(REG2_REG_21__SCAN_IN), .B1(n4293), .B2(
        n4636), .ZN(n4294) );
  OAI21_X1 U4922 ( .B1(n4441), .B2(n4380), .A(n4294), .ZN(n4295) );
  AOI21_X1 U4923 ( .B1(n4296), .B2(n4382), .A(n4295), .ZN(n4297) );
  OAI21_X1 U4924 ( .B1(n4518), .B2(n4385), .A(n4297), .ZN(n4298) );
  AOI21_X1 U4925 ( .B1(n4443), .B2(n4648), .A(n4298), .ZN(n4299) );
  OAI21_X1 U4926 ( .B1(n4300), .B2(n4388), .A(n4299), .ZN(U3269) );
  XNOR2_X1 U4927 ( .A(n4301), .B(n4304), .ZN(n4447) );
  NAND2_X1 U4928 ( .A1(n4303), .A2(n4302), .ZN(n4305) );
  XNOR2_X1 U4929 ( .A(n4305), .B(n4304), .ZN(n4310) );
  AOI22_X1 U4930 ( .A1(n4350), .A2(n4408), .B1(n4306), .B2(n4406), .ZN(n4307)
         );
  OAI21_X1 U4931 ( .B1(n4308), .B2(n4331), .A(n4307), .ZN(n4309) );
  AOI21_X1 U4932 ( .B1(n4310), .B2(n4367), .A(n4309), .ZN(n4311) );
  OAI21_X1 U4933 ( .B1(n4447), .B2(n4312), .A(n4311), .ZN(n4448) );
  NAND2_X1 U4934 ( .A1(n4448), .A2(n4648), .ZN(n4321) );
  INV_X1 U4935 ( .A(n4338), .ZN(n4315) );
  OAI21_X1 U4936 ( .B1(n4315), .B2(n4314), .A(n4313), .ZN(n4522) );
  INV_X1 U4937 ( .A(n4522), .ZN(n4319) );
  INV_X1 U4938 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4317) );
  OAI22_X1 U4939 ( .A1(n4648), .A2(n4317), .B1(n4316), .B2(n4645), .ZN(n4318)
         );
  AOI21_X1 U4940 ( .B1(n4319), .B2(n4652), .A(n4318), .ZN(n4320) );
  OAI211_X1 U4941 ( .C1(n4447), .C2(n4322), .A(n4321), .B(n4320), .ZN(U3270)
         );
  XNOR2_X1 U4942 ( .A(n4323), .B(n4330), .ZN(n4453) );
  INV_X1 U4943 ( .A(n4453), .ZN(n4343) );
  NAND2_X1 U4944 ( .A1(n4325), .A2(n4324), .ZN(n4347) );
  INV_X1 U4945 ( .A(n4326), .ZN(n4328) );
  OAI21_X1 U4946 ( .B1(n4347), .B2(n4328), .A(n4327), .ZN(n4329) );
  XOR2_X1 U4947 ( .A(n4330), .B(n4329), .Z(n4335) );
  OAI22_X1 U4948 ( .A1(n4441), .A2(n4331), .B1(n4459), .B2(n4336), .ZN(n4332)
         );
  AOI21_X1 U4949 ( .B1(n4408), .B2(n4370), .A(n4332), .ZN(n4333) );
  OAI21_X1 U4950 ( .B1(n4335), .B2(n4334), .A(n4333), .ZN(n4452) );
  OR2_X1 U4951 ( .A1(n4355), .A2(n4336), .ZN(n4337) );
  NAND2_X1 U4952 ( .A1(n4338), .A2(n4337), .ZN(n4526) );
  AOI22_X1 U4953 ( .A1(n4378), .A2(REG2_REG_19__SCAN_IN), .B1(n4339), .B2(
        n4636), .ZN(n4340) );
  OAI21_X1 U4954 ( .B1(n4526), .B2(n4385), .A(n4340), .ZN(n4341) );
  AOI21_X1 U4955 ( .B1(n4452), .B2(n4648), .A(n4341), .ZN(n4342) );
  OAI21_X1 U4956 ( .B1(n4343), .B2(n4388), .A(n4342), .ZN(U3271) );
  OAI21_X1 U4957 ( .B1(n4345), .B2(n4348), .A(n4344), .ZN(n4346) );
  INV_X1 U4958 ( .A(n4346), .ZN(n4457) );
  XOR2_X1 U4959 ( .A(n4348), .B(n4347), .Z(n4354) );
  AOI22_X1 U4960 ( .A1(n4350), .A2(n4369), .B1(n4349), .B2(n4406), .ZN(n4351)
         );
  OAI21_X1 U4961 ( .B1(n4352), .B2(n4460), .A(n4351), .ZN(n4353) );
  AOI21_X1 U4962 ( .B1(n4354), .B2(n4367), .A(n4353), .ZN(n4456) );
  INV_X1 U4963 ( .A(n4456), .ZN(n4362) );
  INV_X1 U4964 ( .A(n4355), .ZN(n4356) );
  OAI211_X1 U4965 ( .C1(n4374), .C2(n4357), .A(n4356), .B(n4474), .ZN(n4455)
         );
  AOI22_X1 U4966 ( .A1(n4378), .A2(REG2_REG_18__SCAN_IN), .B1(n4358), .B2(
        n4636), .ZN(n4359) );
  OAI21_X1 U4967 ( .B1(n4455), .B2(n4360), .A(n4359), .ZN(n4361) );
  AOI21_X1 U4968 ( .B1(n4362), .B2(n4648), .A(n4361), .ZN(n4363) );
  OAI21_X1 U4969 ( .B1(n4457), .B2(n4388), .A(n4363), .ZN(U3272) );
  XOR2_X1 U4970 ( .A(n4365), .B(n4364), .Z(n4464) );
  INV_X1 U4971 ( .A(n4464), .ZN(n4389) );
  XNOR2_X1 U4972 ( .A(n4366), .B(n4365), .ZN(n4368) );
  NAND2_X1 U4973 ( .A1(n4368), .A2(n4367), .ZN(n4372) );
  NAND2_X1 U4974 ( .A1(n4370), .A2(n4369), .ZN(n4371) );
  NAND2_X1 U4975 ( .A1(n4372), .A2(n4371), .ZN(n4463) );
  INV_X1 U4976 ( .A(n4373), .ZN(n4376) );
  INV_X1 U4977 ( .A(n4374), .ZN(n4375) );
  OAI21_X1 U4978 ( .B1(n4376), .B2(n4458), .A(n4375), .ZN(n4532) );
  AOI22_X1 U4979 ( .A1(n4378), .A2(REG2_REG_17__SCAN_IN), .B1(n4377), .B2(
        n4636), .ZN(n4379) );
  OAI21_X1 U4980 ( .B1(n4461), .B2(n4380), .A(n4379), .ZN(n4381) );
  AOI21_X1 U4981 ( .B1(n4383), .B2(n4382), .A(n4381), .ZN(n4384) );
  OAI21_X1 U4982 ( .B1(n4532), .B2(n4385), .A(n4384), .ZN(n4386) );
  AOI21_X1 U4983 ( .B1(n4463), .B2(n4648), .A(n4386), .ZN(n4387) );
  OAI21_X1 U4984 ( .B1(n4389), .B2(n4388), .A(n4387), .ZN(U3273) );
  NOR2_X1 U4985 ( .A1(n4713), .A2(n4390), .ZN(n4391) );
  AOI21_X1 U4986 ( .B1(n4713), .B2(n4480), .A(n4391), .ZN(n4392) );
  OAI21_X1 U4987 ( .B1(n4483), .B2(n4467), .A(n4392), .ZN(U3549) );
  AOI21_X1 U4988 ( .B1(n4395), .B2(n4394), .A(n4393), .ZN(n4550) );
  INV_X1 U4989 ( .A(n4550), .ZN(n4486) );
  NAND2_X1 U4990 ( .A1(n4406), .A2(n4395), .ZN(n4396) );
  AND2_X1 U4991 ( .A1(n4397), .A2(n4396), .ZN(n4552) );
  INV_X1 U4992 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4398) );
  MUX2_X1 U4993 ( .A(n4552), .B(n4398), .S(n4710), .Z(n4399) );
  OAI21_X1 U4994 ( .B1(n4486), .B2(n4467), .A(n4399), .ZN(U3548) );
  AOI22_X1 U4995 ( .A1(n4400), .A2(n4408), .B1(n2324), .B2(n4406), .ZN(n4401)
         );
  OAI211_X1 U4996 ( .C1(n4403), .C2(n4468), .A(n4402), .B(n4401), .ZN(n4487)
         );
  MUX2_X1 U4997 ( .A(REG1_REG_28__SCAN_IN), .B(n4487), .S(n4713), .Z(n4404) );
  INV_X1 U4998 ( .A(n4404), .ZN(n4405) );
  OAI21_X1 U4999 ( .B1(n4467), .B2(n4490), .A(n4405), .ZN(U3546) );
  AOI22_X1 U5000 ( .A1(n4409), .A2(n4408), .B1(n4407), .B2(n4406), .ZN(n4410)
         );
  OAI211_X1 U5001 ( .C1(n4412), .C2(n4468), .A(n4411), .B(n4410), .ZN(n4491)
         );
  MUX2_X1 U5002 ( .A(REG1_REG_27__SCAN_IN), .B(n4491), .S(n4713), .Z(n4413) );
  INV_X1 U5003 ( .A(n4413), .ZN(n4414) );
  OAI21_X1 U5004 ( .B1(n4467), .B2(n4494), .A(n4414), .ZN(U3545) );
  INV_X1 U5005 ( .A(n4415), .ZN(n4416) );
  AOI21_X1 U5006 ( .B1(n4417), .B2(n4688), .A(n4416), .ZN(n4495) );
  MUX2_X1 U5007 ( .A(n4418), .B(n4495), .S(n4713), .Z(n4419) );
  OAI21_X1 U5008 ( .B1(n4467), .B2(n4498), .A(n4419), .ZN(U3544) );
  AOI21_X1 U5009 ( .B1(n4421), .B2(n4688), .A(n4420), .ZN(n4499) );
  MUX2_X1 U5010 ( .A(n4422), .B(n4499), .S(n4713), .Z(n4423) );
  OAI21_X1 U5011 ( .B1(n4467), .B2(n4502), .A(n4423), .ZN(U3543) );
  INV_X1 U5012 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4429) );
  OAI22_X1 U5013 ( .A1(n4425), .A2(n4460), .B1(n4424), .B2(n4459), .ZN(n4426)
         );
  AOI211_X1 U5014 ( .C1(n4428), .C2(n4688), .A(n4427), .B(n4426), .ZN(n4503)
         );
  MUX2_X1 U5015 ( .A(n4429), .B(n4503), .S(n4713), .Z(n4430) );
  OAI21_X1 U5016 ( .B1(n4467), .B2(n4506), .A(n4430), .ZN(U3542) );
  AOI21_X1 U5017 ( .B1(n4432), .B2(n4688), .A(n4431), .ZN(n4507) );
  MUX2_X1 U5018 ( .A(n4433), .B(n4507), .S(n4713), .Z(n4434) );
  OAI21_X1 U5019 ( .B1(n4467), .B2(n4510), .A(n4434), .ZN(U3541) );
  INV_X1 U5020 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4438) );
  INV_X1 U5021 ( .A(n4435), .ZN(n4437) );
  AOI21_X1 U5022 ( .B1(n4437), .B2(n4688), .A(n4436), .ZN(n4511) );
  MUX2_X1 U5023 ( .A(n4438), .B(n4511), .S(n4713), .Z(n4439) );
  OAI21_X1 U5024 ( .B1(n4467), .B2(n4514), .A(n4439), .ZN(U3540) );
  INV_X1 U5025 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4445) );
  OAI22_X1 U5026 ( .A1(n4441), .A2(n4460), .B1(n4459), .B2(n4440), .ZN(n4442)
         );
  AOI211_X1 U5027 ( .C1(n4444), .C2(n4688), .A(n4443), .B(n4442), .ZN(n4515)
         );
  MUX2_X1 U5028 ( .A(n4445), .B(n4515), .S(n4713), .Z(n4446) );
  OAI21_X1 U5029 ( .B1(n4467), .B2(n4518), .A(n4446), .ZN(U3539) );
  INV_X1 U5030 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4450) );
  INV_X1 U5031 ( .A(n4447), .ZN(n4449) );
  AOI21_X1 U5032 ( .B1(n4699), .B2(n4449), .A(n4448), .ZN(n4519) );
  MUX2_X1 U5033 ( .A(n4450), .B(n4519), .S(n4713), .Z(n4451) );
  OAI21_X1 U5034 ( .B1(n4467), .B2(n4522), .A(n4451), .ZN(U3538) );
  AOI21_X1 U5035 ( .B1(n4453), .B2(n4688), .A(n4452), .ZN(n4523) );
  MUX2_X1 U5036 ( .A(n4137), .B(n4523), .S(n4713), .Z(n4454) );
  OAI21_X1 U5037 ( .B1(n4467), .B2(n4526), .A(n4454), .ZN(U3537) );
  OAI211_X1 U5038 ( .C1(n4457), .C2(n4468), .A(n4456), .B(n4455), .ZN(n4527)
         );
  MUX2_X1 U5039 ( .A(REG1_REG_18__SCAN_IN), .B(n4527), .S(n4713), .Z(U3536) );
  INV_X1 U5040 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4465) );
  OAI22_X1 U5041 ( .A1(n4461), .A2(n4460), .B1(n4459), .B2(n4458), .ZN(n4462)
         );
  AOI211_X1 U5042 ( .C1(n4464), .C2(n4688), .A(n4463), .B(n4462), .ZN(n4528)
         );
  MUX2_X1 U5043 ( .A(n4465), .B(n4528), .S(n4713), .Z(n4466) );
  OAI21_X1 U5044 ( .B1(n4467), .B2(n4532), .A(n4466), .ZN(U3535) );
  OR2_X1 U5045 ( .A1(n4469), .A2(n4468), .ZN(n4471) );
  NAND2_X1 U5046 ( .A1(n4471), .A2(n4470), .ZN(n4533) );
  MUX2_X1 U5047 ( .A(n4533), .B(REG1_REG_16__SCAN_IN), .S(n4710), .Z(n4473) );
  NOR2_X1 U5048 ( .A1(n4534), .A2(n4467), .ZN(n4472) );
  NAND3_X1 U5049 ( .A1(n4476), .A2(n4475), .A3(n4474), .ZN(n4477) );
  OAI211_X1 U5050 ( .C1(n4479), .C2(n4674), .A(n4478), .B(n4477), .ZN(n4537)
         );
  MUX2_X1 U5051 ( .A(REG1_REG_14__SCAN_IN), .B(n4537), .S(n4713), .Z(U3532) );
  NAND2_X1 U5052 ( .A1(n4702), .A2(n4480), .ZN(n4482) );
  NAND2_X1 U5053 ( .A1(n4700), .A2(REG0_REG_31__SCAN_IN), .ZN(n4481) );
  OAI211_X1 U5054 ( .C1(n4483), .C2(n4531), .A(n4482), .B(n4481), .ZN(U3517)
         );
  INV_X1 U5055 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4484) );
  MUX2_X1 U5056 ( .A(n4552), .B(n4484), .S(n4700), .Z(n4485) );
  OAI21_X1 U5057 ( .B1(n4486), .B2(n4531), .A(n4485), .ZN(U3516) );
  MUX2_X1 U5058 ( .A(REG0_REG_28__SCAN_IN), .B(n4487), .S(n4702), .Z(n4488) );
  INV_X1 U5059 ( .A(n4488), .ZN(n4489) );
  OAI21_X1 U5060 ( .B1(n4490), .B2(n4531), .A(n4489), .ZN(U3514) );
  MUX2_X1 U5061 ( .A(REG0_REG_27__SCAN_IN), .B(n4491), .S(n4702), .Z(n4492) );
  INV_X1 U5062 ( .A(n4492), .ZN(n4493) );
  OAI21_X1 U5063 ( .B1(n4494), .B2(n4531), .A(n4493), .ZN(U3513) );
  INV_X1 U5064 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4496) );
  MUX2_X1 U5065 ( .A(n4496), .B(n4495), .S(n4702), .Z(n4497) );
  OAI21_X1 U5066 ( .B1(n4498), .B2(n4531), .A(n4497), .ZN(U3512) );
  INV_X1 U5067 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4500) );
  MUX2_X1 U5068 ( .A(n4500), .B(n4499), .S(n4702), .Z(n4501) );
  OAI21_X1 U5069 ( .B1(n4502), .B2(n4531), .A(n4501), .ZN(U3511) );
  INV_X1 U5070 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4504) );
  MUX2_X1 U5071 ( .A(n4504), .B(n4503), .S(n4702), .Z(n4505) );
  OAI21_X1 U5072 ( .B1(n4506), .B2(n4531), .A(n4505), .ZN(U3510) );
  INV_X1 U5073 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4508) );
  MUX2_X1 U5074 ( .A(n4508), .B(n4507), .S(n4702), .Z(n4509) );
  OAI21_X1 U5075 ( .B1(n4510), .B2(n4531), .A(n4509), .ZN(U3509) );
  INV_X1 U5076 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4512) );
  MUX2_X1 U5077 ( .A(n4512), .B(n4511), .S(n4702), .Z(n4513) );
  OAI21_X1 U5078 ( .B1(n4514), .B2(n4531), .A(n4513), .ZN(U3508) );
  INV_X1 U5079 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4516) );
  MUX2_X1 U5080 ( .A(n4516), .B(n4515), .S(n4702), .Z(n4517) );
  OAI21_X1 U5081 ( .B1(n4518), .B2(n4531), .A(n4517), .ZN(U3507) );
  INV_X1 U5082 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4520) );
  MUX2_X1 U5083 ( .A(n4520), .B(n4519), .S(n4702), .Z(n4521) );
  OAI21_X1 U5084 ( .B1(n4522), .B2(n4531), .A(n4521), .ZN(U3506) );
  INV_X1 U5085 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4524) );
  MUX2_X1 U5086 ( .A(n4524), .B(n4523), .S(n4702), .Z(n4525) );
  OAI21_X1 U5087 ( .B1(n4526), .B2(n4531), .A(n4525), .ZN(U3505) );
  MUX2_X1 U5088 ( .A(REG0_REG_18__SCAN_IN), .B(n4527), .S(n4702), .Z(U3503) );
  INV_X1 U5089 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4529) );
  MUX2_X1 U5090 ( .A(n4529), .B(n4528), .S(n4702), .Z(n4530) );
  OAI21_X1 U5091 ( .B1(n4532), .B2(n4531), .A(n4530), .ZN(U3501) );
  MUX2_X1 U5092 ( .A(n4533), .B(REG0_REG_16__SCAN_IN), .S(n4700), .Z(n4536) );
  NOR2_X1 U5093 ( .A1(n4534), .A2(n4531), .ZN(n4535) );
  MUX2_X1 U5094 ( .A(REG0_REG_14__SCAN_IN), .B(n4537), .S(n4702), .Z(U3495) );
  MUX2_X1 U5095 ( .A(n4538), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5096 ( .A(n4539), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5097 ( .A(n4540), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5098 ( .A(n4541), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U5099 ( .A(n4553), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5100 ( .A(DATAI_8_), .B(n4542), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5101 ( .A(n4543), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5102 ( .A(n4544), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5103 ( .A(n4545), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5104 ( .A(DATAI_4_), .B(n4546), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5105 ( .A(n4547), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5106 ( .A(n4548), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5107 ( .A(n4549), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U5108 ( .A1(n4550), .A2(n4652), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4378), .ZN(n4551) );
  OAI21_X1 U5109 ( .B1(n4378), .B2(n4552), .A(n4551), .ZN(U3261) );
  INV_X1 U5110 ( .A(n4553), .ZN(n4562) );
  OAI211_X1 U5111 ( .C1(n4556), .C2(n4555), .A(n4587), .B(n4554), .ZN(n4561)
         );
  OAI211_X1 U5112 ( .C1(n4559), .C2(n4558), .A(n4629), .B(n4557), .ZN(n4560)
         );
  OAI211_X1 U5113 ( .C1(n4635), .C2(n4562), .A(n4561), .B(n4560), .ZN(n4563)
         );
  AOI211_X1 U5114 ( .C1(n4628), .C2(ADDR_REG_9__SCAN_IN), .A(n4564), .B(n4563), 
        .ZN(n4565) );
  INV_X1 U5115 ( .A(n4565), .ZN(U3249) );
  OAI211_X1 U5116 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4567), .A(n4587), .B(n4566), .ZN(n4569) );
  NAND2_X1 U5117 ( .A1(n4569), .A2(n4568), .ZN(n4570) );
  AOI21_X1 U5118 ( .B1(n4628), .B2(ADDR_REG_10__SCAN_IN), .A(n4570), .ZN(n4574) );
  OAI211_X1 U5119 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4572), .A(n4629), .B(n4571), .ZN(n4573) );
  OAI211_X1 U5120 ( .C1(n4635), .C2(n4668), .A(n4574), .B(n4573), .ZN(U3250)
         );
  OAI211_X1 U5121 ( .C1(n4577), .C2(n4576), .A(n4629), .B(n4575), .ZN(n4582)
         );
  OAI211_X1 U5122 ( .C1(n4580), .C2(n4579), .A(n4587), .B(n4578), .ZN(n4581)
         );
  OAI211_X1 U5123 ( .C1(n4635), .C2(n4667), .A(n4582), .B(n4581), .ZN(n4583)
         );
  AOI211_X1 U5124 ( .C1(n4628), .C2(ADDR_REG_11__SCAN_IN), .A(n4584), .B(n4583), .ZN(n4585) );
  INV_X1 U5125 ( .A(n4585), .ZN(U3251) );
  OAI211_X1 U5126 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4588), .A(n4587), .B(n4586), .ZN(n4590) );
  NAND2_X1 U5127 ( .A1(n4590), .A2(n4589), .ZN(n4591) );
  AOI21_X1 U5128 ( .B1(n4628), .B2(ADDR_REG_12__SCAN_IN), .A(n4591), .ZN(n4595) );
  OAI211_X1 U5129 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4593), .A(n4629), .B(n4592), .ZN(n4594) );
  OAI211_X1 U5130 ( .C1(n4635), .C2(n4665), .A(n4595), .B(n4594), .ZN(U3252)
         );
  AOI211_X1 U5131 ( .C1(n4598), .C2(n4597), .A(n4596), .B(n4622), .ZN(n4599)
         );
  AOI211_X1 U5132 ( .C1(n4628), .C2(ADDR_REG_14__SCAN_IN), .A(n4600), .B(n4599), .ZN(n4604) );
  OAI211_X1 U5133 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4602), .A(n4629), .B(n4601), .ZN(n4603) );
  OAI211_X1 U5134 ( .C1(n4635), .C2(n2336), .A(n4604), .B(n4603), .ZN(U3254)
         );
  AOI211_X1 U5135 ( .C1(n4606), .C2(n4605), .A(n2248), .B(n4622), .ZN(n4607)
         );
  AOI211_X1 U5136 ( .C1(n4628), .C2(ADDR_REG_15__SCAN_IN), .A(n4608), .B(n4607), .ZN(n4613) );
  OAI211_X1 U5137 ( .C1(n4611), .C2(n4610), .A(n4629), .B(n4609), .ZN(n4612)
         );
  OAI211_X1 U5138 ( .C1(n4635), .C2(n4664), .A(n4613), .B(n4612), .ZN(U3255)
         );
  AOI221_X1 U5139 ( .B1(n4615), .B2(n4614), .C1(n3610), .C2(n4614), .A(n4622), 
        .ZN(n4616) );
  AOI211_X1 U5140 ( .C1(n4628), .C2(ADDR_REG_16__SCAN_IN), .A(n4617), .B(n4616), .ZN(n4621) );
  OAI221_X1 U5141 ( .B1(n4619), .B2(REG1_REG_16__SCAN_IN), .C1(n4619), .C2(
        n4618), .A(n4629), .ZN(n4620) );
  OAI211_X1 U5142 ( .C1(n4635), .C2(n4663), .A(n4621), .B(n4620), .ZN(U3256)
         );
  AOI221_X1 U5143 ( .B1(n4625), .B2(n4624), .C1(n4623), .C2(n4624), .A(n4622), 
        .ZN(n4626) );
  AOI211_X1 U5144 ( .C1(n4628), .C2(ADDR_REG_17__SCAN_IN), .A(n4627), .B(n4626), .ZN(n4634) );
  OAI221_X1 U5145 ( .B1(n4632), .B2(n4631), .C1(n4632), .C2(n4630), .A(n4629), 
        .ZN(n4633) );
  OAI211_X1 U5146 ( .C1(n4635), .C2(n4662), .A(n4634), .B(n4633), .ZN(U3257)
         );
  AOI22_X1 U5147 ( .A1(n4637), .A2(n4636), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4378), .ZN(n4642) );
  INV_X1 U5148 ( .A(n4638), .ZN(n4639) );
  AOI22_X1 U5149 ( .A1(n4640), .A2(n4653), .B1(n4652), .B2(n4639), .ZN(n4641)
         );
  OAI211_X1 U5150 ( .C1(n4378), .C2(n4643), .A(n4642), .B(n4641), .ZN(U3280)
         );
  INV_X1 U5151 ( .A(n4644), .ZN(n4646) );
  OAI22_X1 U5152 ( .A1(n4648), .A2(n4647), .B1(n4646), .B2(n4645), .ZN(n4649)
         );
  INV_X1 U5153 ( .A(n4649), .ZN(n4656) );
  INV_X1 U5154 ( .A(n4650), .ZN(n4651) );
  AOI22_X1 U5155 ( .A1(n4654), .A2(n4653), .B1(n4652), .B2(n4651), .ZN(n4655)
         );
  OAI211_X1 U5156 ( .C1(n4378), .C2(n4657), .A(n4656), .B(n4655), .ZN(U3282)
         );
  AND2_X1 U5157 ( .A1(n4659), .A2(D_REG_31__SCAN_IN), .ZN(U3291) );
  INV_X1 U5158 ( .A(D_REG_30__SCAN_IN), .ZN(n4855) );
  NOR2_X1 U5159 ( .A1(n4658), .A2(n4855), .ZN(U3292) );
  INV_X1 U5160 ( .A(D_REG_29__SCAN_IN), .ZN(n5054) );
  NOR2_X1 U5161 ( .A1(n4658), .A2(n5054), .ZN(U3293) );
  INV_X1 U5162 ( .A(D_REG_28__SCAN_IN), .ZN(n5092) );
  NOR2_X1 U5163 ( .A1(n4658), .A2(n5092), .ZN(U3294) );
  AND2_X1 U5164 ( .A1(n4659), .A2(D_REG_27__SCAN_IN), .ZN(U3295) );
  INV_X1 U5165 ( .A(D_REG_26__SCAN_IN), .ZN(n4880) );
  NOR2_X1 U5166 ( .A1(n4658), .A2(n4880), .ZN(U3296) );
  INV_X1 U5167 ( .A(D_REG_25__SCAN_IN), .ZN(n4812) );
  NOR2_X1 U5168 ( .A1(n4658), .A2(n4812), .ZN(U3297) );
  INV_X1 U5169 ( .A(D_REG_24__SCAN_IN), .ZN(n4881) );
  NOR2_X1 U5170 ( .A1(n4658), .A2(n4881), .ZN(U3298) );
  INV_X1 U5171 ( .A(D_REG_23__SCAN_IN), .ZN(n5046) );
  NOR2_X1 U5172 ( .A1(n4658), .A2(n5046), .ZN(U3299) );
  INV_X1 U5173 ( .A(D_REG_22__SCAN_IN), .ZN(n5043) );
  NOR2_X1 U5174 ( .A1(n4658), .A2(n5043), .ZN(U3300) );
  INV_X1 U5175 ( .A(D_REG_21__SCAN_IN), .ZN(n4871) );
  NOR2_X1 U5176 ( .A1(n4658), .A2(n4871), .ZN(U3301) );
  INV_X1 U5177 ( .A(D_REG_20__SCAN_IN), .ZN(n5047) );
  NOR2_X1 U5178 ( .A1(n4658), .A2(n5047), .ZN(U3302) );
  INV_X1 U5179 ( .A(D_REG_19__SCAN_IN), .ZN(n4841) );
  NOR2_X1 U5180 ( .A1(n4658), .A2(n4841), .ZN(U3303) );
  INV_X1 U5181 ( .A(D_REG_18__SCAN_IN), .ZN(n5040) );
  NOR2_X1 U5182 ( .A1(n4658), .A2(n5040), .ZN(U3304) );
  INV_X1 U5183 ( .A(D_REG_17__SCAN_IN), .ZN(n5044) );
  NOR2_X1 U5184 ( .A1(n4658), .A2(n5044), .ZN(U3305) );
  INV_X1 U5185 ( .A(D_REG_16__SCAN_IN), .ZN(n4786) );
  NOR2_X1 U5186 ( .A1(n4658), .A2(n4786), .ZN(U3306) );
  INV_X1 U5187 ( .A(D_REG_15__SCAN_IN), .ZN(n5059) );
  NOR2_X1 U5188 ( .A1(n4658), .A2(n5059), .ZN(U3307) );
  AND2_X1 U5189 ( .A1(n4659), .A2(D_REG_14__SCAN_IN), .ZN(U3308) );
  AND2_X1 U5190 ( .A1(n4659), .A2(D_REG_13__SCAN_IN), .ZN(U3309) );
  INV_X1 U5191 ( .A(D_REG_12__SCAN_IN), .ZN(n4808) );
  NOR2_X1 U5192 ( .A1(n4658), .A2(n4808), .ZN(U3310) );
  INV_X1 U5193 ( .A(D_REG_11__SCAN_IN), .ZN(n4815) );
  NOR2_X1 U5194 ( .A1(n4658), .A2(n4815), .ZN(U3311) );
  INV_X1 U5195 ( .A(D_REG_10__SCAN_IN), .ZN(n4847) );
  NOR2_X1 U5196 ( .A1(n4658), .A2(n4847), .ZN(U3312) );
  INV_X1 U5197 ( .A(D_REG_9__SCAN_IN), .ZN(n5041) );
  NOR2_X1 U5198 ( .A1(n4658), .A2(n5041), .ZN(U3313) );
  INV_X1 U5199 ( .A(D_REG_8__SCAN_IN), .ZN(n5038) );
  NOR2_X1 U5200 ( .A1(n4658), .A2(n5038), .ZN(U3314) );
  INV_X1 U5201 ( .A(D_REG_7__SCAN_IN), .ZN(n5056) );
  NOR2_X1 U5202 ( .A1(n4658), .A2(n5056), .ZN(U3315) );
  INV_X1 U5203 ( .A(D_REG_6__SCAN_IN), .ZN(n5053) );
  NOR2_X1 U5204 ( .A1(n4658), .A2(n5053), .ZN(U3316) );
  INV_X1 U5205 ( .A(D_REG_5__SCAN_IN), .ZN(n4764) );
  NOR2_X1 U5206 ( .A1(n4658), .A2(n4764), .ZN(U3317) );
  INV_X1 U5207 ( .A(D_REG_4__SCAN_IN), .ZN(n5060) );
  NOR2_X1 U5208 ( .A1(n4658), .A2(n5060), .ZN(U3318) );
  INV_X1 U5209 ( .A(D_REG_3__SCAN_IN), .ZN(n5057) );
  NOR2_X1 U5210 ( .A1(n4658), .A2(n5057), .ZN(U3319) );
  AND2_X1 U5211 ( .A1(n4659), .A2(D_REG_2__SCAN_IN), .ZN(U3320) );
  INV_X1 U5212 ( .A(DATAI_23_), .ZN(n4978) );
  AOI21_X1 U5213 ( .B1(U3149), .B2(n4978), .A(n4660), .ZN(U3329) );
  AOI22_X1 U5214 ( .A1(STATE_REG_SCAN_IN), .A2(n4662), .B1(n4661), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5215 ( .A(DATAI_16_), .ZN(n4867) );
  AOI22_X1 U5216 ( .A1(STATE_REG_SCAN_IN), .A2(n4663), .B1(n4867), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5217 ( .A(DATAI_15_), .ZN(n4983) );
  AOI22_X1 U5218 ( .A1(STATE_REG_SCAN_IN), .A2(n4664), .B1(n4983), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5219 ( .A(DATAI_14_), .ZN(n4995) );
  AOI22_X1 U5220 ( .A1(STATE_REG_SCAN_IN), .A2(n2336), .B1(n4995), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5221 ( .A(DATAI_12_), .ZN(n4816) );
  AOI22_X1 U5222 ( .A1(STATE_REG_SCAN_IN), .A2(n4665), .B1(n4816), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5223 ( .A(DATAI_11_), .ZN(n4666) );
  AOI22_X1 U5224 ( .A1(STATE_REG_SCAN_IN), .A2(n4667), .B1(n4666), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5225 ( .A(DATAI_10_), .ZN(n4828) );
  AOI22_X1 U5226 ( .A1(STATE_REG_SCAN_IN), .A2(n4668), .B1(n4828), .B2(U3149), 
        .ZN(U3342) );
  OAI211_X1 U5227 ( .C1(n4671), .C2(n4674), .A(n4670), .B(n4669), .ZN(n4672)
         );
  INV_X1 U5228 ( .A(n4672), .ZN(n4703) );
  INV_X1 U5229 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4856) );
  AOI22_X1 U5230 ( .A1(n4702), .A2(n4703), .B1(n4856), .B2(n4700), .ZN(U3467)
         );
  OAI22_X1 U5231 ( .A1(n4675), .A2(n4674), .B1(n4694), .B2(n4673), .ZN(n4676)
         );
  NOR2_X1 U5232 ( .A1(n4677), .A2(n4676), .ZN(n4704) );
  INV_X1 U5233 ( .A(REG0_REG_1__SCAN_IN), .ZN(n5026) );
  AOI22_X1 U5234 ( .A1(n4702), .A2(n4704), .B1(n5026), .B2(n4700), .ZN(U3469)
         );
  NOR3_X1 U5235 ( .A1(n4679), .A2(n4678), .A3(n4694), .ZN(n4681) );
  AOI211_X1 U5236 ( .C1(n4699), .C2(n4682), .A(n4681), .B(n4680), .ZN(n4705)
         );
  INV_X1 U5237 ( .A(REG0_REG_2__SCAN_IN), .ZN(n5061) );
  AOI22_X1 U5238 ( .A1(n4702), .A2(n4705), .B1(n5061), .B2(n4700), .ZN(U3471)
         );
  INV_X1 U5239 ( .A(n4683), .ZN(n4685) );
  AOI211_X1 U5240 ( .C1(n4686), .C2(n4699), .A(n4685), .B(n4684), .ZN(n4707)
         );
  INV_X1 U5241 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4687) );
  AOI22_X1 U5242 ( .A1(n4702), .A2(n4707), .B1(n4687), .B2(n4700), .ZN(U3475)
         );
  NAND2_X1 U5243 ( .A1(n4689), .A2(n4688), .ZN(n4691) );
  INV_X1 U5244 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4693) );
  AOI22_X1 U5245 ( .A1(n4702), .A2(n4709), .B1(n4693), .B2(n4700), .ZN(U3481)
         );
  NOR2_X1 U5246 ( .A1(n4695), .A2(n4694), .ZN(n4697) );
  AOI211_X1 U5247 ( .C1(n4699), .C2(n4698), .A(n4697), .B(n4696), .ZN(n4712)
         );
  INV_X1 U5248 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4701) );
  AOI22_X1 U5249 ( .A1(n4702), .A2(n4712), .B1(n4701), .B2(n4700), .ZN(U3489)
         );
  AOI22_X1 U5250 ( .A1(n4713), .A2(n4703), .B1(n2530), .B2(n4710), .ZN(U3518)
         );
  AOI22_X1 U5251 ( .A1(n4713), .A2(n4704), .B1(n2545), .B2(n4710), .ZN(U3519)
         );
  AOI22_X1 U5252 ( .A1(n4713), .A2(n4705), .B1(n2563), .B2(n4710), .ZN(U3520)
         );
  INV_X1 U5253 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4706) );
  AOI22_X1 U5254 ( .A1(n4713), .A2(n4707), .B1(n4706), .B2(n4710), .ZN(U3522)
         );
  AOI22_X1 U5255 ( .A1(n4713), .A2(n4709), .B1(n4708), .B2(n4710), .ZN(U3525)
         );
  AOI22_X1 U5256 ( .A1(n4713), .A2(n4712), .B1(n4711), .B2(n4710), .ZN(U3529)
         );
  OAI22_X1 U5257 ( .A1(DATAI_25_), .A2(keyinput_g6), .B1(DATAI_24_), .B2(
        keyinput_g7), .ZN(n4714) );
  AOI221_X1 U5258 ( .B1(DATAI_25_), .B2(keyinput_g6), .C1(keyinput_g7), .C2(
        DATAI_24_), .A(n4714), .ZN(n4721) );
  OAI22_X1 U5259 ( .A1(IR_REG_28__SCAN_IN), .A2(keyinput_g83), .B1(
        keyinput_g126), .B2(REG0_REG_7__SCAN_IN), .ZN(n4715) );
  AOI221_X1 U5260 ( .B1(IR_REG_28__SCAN_IN), .B2(keyinput_g83), .C1(
        REG0_REG_7__SCAN_IN), .C2(keyinput_g126), .A(n4715), .ZN(n4720) );
  OAI22_X1 U5261 ( .A1(DATAI_14_), .A2(keyinput_g17), .B1(REG0_REG_1__SCAN_IN), 
        .B2(keyinput_g120), .ZN(n4716) );
  AOI221_X1 U5262 ( .B1(DATAI_14_), .B2(keyinput_g17), .C1(keyinput_g120), 
        .C2(REG0_REG_1__SCAN_IN), .A(n4716), .ZN(n4719) );
  OAI22_X1 U5263 ( .A1(IR_REG_20__SCAN_IN), .A2(keyinput_g75), .B1(
        D_REG_23__SCAN_IN), .B2(keyinput_g110), .ZN(n4717) );
  AOI221_X1 U5264 ( .B1(IR_REG_20__SCAN_IN), .B2(keyinput_g75), .C1(
        keyinput_g110), .C2(D_REG_23__SCAN_IN), .A(n4717), .ZN(n4718) );
  NAND4_X1 U5265 ( .A1(n4721), .A2(n4720), .A3(n4719), .A4(n4718), .ZN(n4749)
         );
  OAI22_X1 U5266 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput_g46), .B1(DATAI_17_), .B2(keyinput_g14), .ZN(n4722) );
  AOI221_X1 U5267 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput_g46), .C1(
        keyinput_g14), .C2(DATAI_17_), .A(n4722), .ZN(n4729) );
  OAI22_X1 U5268 ( .A1(IR_REG_15__SCAN_IN), .A2(keyinput_g70), .B1(
        keyinput_g100), .B2(D_REG_13__SCAN_IN), .ZN(n4723) );
  AOI221_X1 U5269 ( .B1(IR_REG_15__SCAN_IN), .B2(keyinput_g70), .C1(
        D_REG_13__SCAN_IN), .C2(keyinput_g100), .A(n4723), .ZN(n4728) );
  OAI22_X1 U5270 ( .A1(IR_REG_12__SCAN_IN), .A2(keyinput_g67), .B1(
        keyinput_g124), .B2(REG0_REG_5__SCAN_IN), .ZN(n4724) );
  AOI221_X1 U5271 ( .B1(IR_REG_12__SCAN_IN), .B2(keyinput_g67), .C1(
        REG0_REG_5__SCAN_IN), .C2(keyinput_g124), .A(n4724), .ZN(n4727) );
  OAI22_X1 U5272 ( .A1(D_REG_9__SCAN_IN), .A2(keyinput_g96), .B1(keyinput_g30), 
        .B2(DATAI_1_), .ZN(n4725) );
  AOI221_X1 U5273 ( .B1(D_REG_9__SCAN_IN), .B2(keyinput_g96), .C1(DATAI_1_), 
        .C2(keyinput_g30), .A(n4725), .ZN(n4726) );
  NAND4_X1 U5274 ( .A1(n4729), .A2(n4728), .A3(n4727), .A4(n4726), .ZN(n4748)
         );
  OAI22_X1 U5275 ( .A1(D_REG_3__SCAN_IN), .A2(keyinput_g90), .B1(DATAI_26_), 
        .B2(keyinput_g5), .ZN(n4730) );
  AOI221_X1 U5276 ( .B1(D_REG_3__SCAN_IN), .B2(keyinput_g90), .C1(keyinput_g5), 
        .C2(DATAI_26_), .A(n4730), .ZN(n4737) );
  OAI22_X1 U5277 ( .A1(DATAI_0_), .A2(keyinput_g31), .B1(keyinput_g123), .B2(
        REG0_REG_4__SCAN_IN), .ZN(n4731) );
  AOI221_X1 U5278 ( .B1(DATAI_0_), .B2(keyinput_g31), .C1(REG0_REG_4__SCAN_IN), 
        .C2(keyinput_g123), .A(n4731), .ZN(n4736) );
  OAI22_X1 U5279 ( .A1(D_REG_18__SCAN_IN), .A2(keyinput_g105), .B1(
        D_REG_17__SCAN_IN), .B2(keyinput_g104), .ZN(n4732) );
  AOI221_X1 U5280 ( .B1(D_REG_18__SCAN_IN), .B2(keyinput_g105), .C1(
        keyinput_g104), .C2(D_REG_17__SCAN_IN), .A(n4732), .ZN(n4735) );
  OAI22_X1 U5281 ( .A1(IR_REG_26__SCAN_IN), .A2(keyinput_g81), .B1(
        REG3_REG_23__SCAN_IN), .B2(keyinput_g36), .ZN(n4733) );
  AOI221_X1 U5282 ( .B1(IR_REG_26__SCAN_IN), .B2(keyinput_g81), .C1(
        keyinput_g36), .C2(REG3_REG_23__SCAN_IN), .A(n4733), .ZN(n4734) );
  NAND4_X1 U5283 ( .A1(n4737), .A2(n4736), .A3(n4735), .A4(n4734), .ZN(n4747)
         );
  OAI22_X1 U5284 ( .A1(IR_REG_24__SCAN_IN), .A2(keyinput_g79), .B1(
        STATE_REG_SCAN_IN), .B2(keyinput_g32), .ZN(n4738) );
  AOI221_X1 U5285 ( .B1(IR_REG_24__SCAN_IN), .B2(keyinput_g79), .C1(
        keyinput_g32), .C2(STATE_REG_SCAN_IN), .A(n4738), .ZN(n4745) );
  OAI22_X1 U5286 ( .A1(REG3_REG_13__SCAN_IN), .A2(keyinput_g54), .B1(
        keyinput_g33), .B2(REG3_REG_7__SCAN_IN), .ZN(n4739) );
  AOI221_X1 U5287 ( .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_g54), .C1(
        REG3_REG_7__SCAN_IN), .C2(keyinput_g33), .A(n4739), .ZN(n4744) );
  OAI22_X1 U5288 ( .A1(D_REG_2__SCAN_IN), .A2(keyinput_g89), .B1(keyinput_g35), 
        .B2(REG3_REG_14__SCAN_IN), .ZN(n4740) );
  AOI221_X1 U5289 ( .B1(D_REG_2__SCAN_IN), .B2(keyinput_g89), .C1(
        REG3_REG_14__SCAN_IN), .C2(keyinput_g35), .A(n4740), .ZN(n4743) );
  OAI22_X1 U5290 ( .A1(REG3_REG_12__SCAN_IN), .A2(keyinput_g44), .B1(
        keyinput_g24), .B2(DATAI_7_), .ZN(n4741) );
  AOI221_X1 U5291 ( .B1(REG3_REG_12__SCAN_IN), .B2(keyinput_g44), .C1(DATAI_7_), .C2(keyinput_g24), .A(n4741), .ZN(n4742) );
  NAND4_X1 U5292 ( .A1(n4745), .A2(n4744), .A3(n4743), .A4(n4742), .ZN(n4746)
         );
  NOR4_X1 U5293 ( .A1(n4749), .A2(n4748), .A3(n4747), .A4(n4746), .ZN(n5097)
         );
  OAI22_X1 U5294 ( .A1(IR_REG_23__SCAN_IN), .A2(keyinput_g78), .B1(
        keyinput_g22), .B2(DATAI_9_), .ZN(n4750) );
  AOI221_X1 U5295 ( .B1(IR_REG_23__SCAN_IN), .B2(keyinput_g78), .C1(DATAI_9_), 
        .C2(keyinput_g22), .A(n4750), .ZN(n4757) );
  OAI22_X1 U5296 ( .A1(REG3_REG_20__SCAN_IN), .A2(keyinput_g53), .B1(
        keyinput_g52), .B2(REG3_REG_0__SCAN_IN), .ZN(n4751) );
  AOI221_X1 U5297 ( .B1(REG3_REG_20__SCAN_IN), .B2(keyinput_g53), .C1(
        REG3_REG_0__SCAN_IN), .C2(keyinput_g52), .A(n4751), .ZN(n4756) );
  OAI22_X1 U5298 ( .A1(DATAI_28_), .A2(keyinput_g3), .B1(keyinput_g1), .B2(
        DATAI_30_), .ZN(n4752) );
  AOI221_X1 U5299 ( .B1(DATAI_28_), .B2(keyinput_g3), .C1(DATAI_30_), .C2(
        keyinput_g1), .A(n4752), .ZN(n4755) );
  OAI22_X1 U5300 ( .A1(DATAI_21_), .A2(keyinput_g10), .B1(DATAI_20_), .B2(
        keyinput_g11), .ZN(n4753) );
  AOI221_X1 U5301 ( .B1(DATAI_21_), .B2(keyinput_g10), .C1(keyinput_g11), .C2(
        DATAI_20_), .A(n4753), .ZN(n4754) );
  NAND4_X1 U5302 ( .A1(n4757), .A2(n4756), .A3(n4755), .A4(n4754), .ZN(n4899)
         );
  OAI22_X1 U5303 ( .A1(DATAI_19_), .A2(keyinput_g12), .B1(DATAI_15_), .B2(
        keyinput_g16), .ZN(n4758) );
  AOI221_X1 U5304 ( .B1(DATAI_19_), .B2(keyinput_g12), .C1(keyinput_g16), .C2(
        DATAI_15_), .A(n4758), .ZN(n4784) );
  OAI22_X1 U5305 ( .A1(D_REG_20__SCAN_IN), .A2(keyinput_g107), .B1(
        D_REG_6__SCAN_IN), .B2(keyinput_g93), .ZN(n4759) );
  AOI221_X1 U5306 ( .B1(D_REG_20__SCAN_IN), .B2(keyinput_g107), .C1(
        keyinput_g93), .C2(D_REG_6__SCAN_IN), .A(n4759), .ZN(n4762) );
  OAI22_X1 U5307 ( .A1(D_REG_27__SCAN_IN), .A2(keyinput_g114), .B1(
        D_REG_22__SCAN_IN), .B2(keyinput_g109), .ZN(n4760) );
  AOI221_X1 U5308 ( .B1(D_REG_27__SCAN_IN), .B2(keyinput_g114), .C1(
        keyinput_g109), .C2(D_REG_22__SCAN_IN), .A(n4760), .ZN(n4761) );
  OAI211_X1 U5309 ( .C1(n4764), .C2(keyinput_g92), .A(n4762), .B(n4761), .ZN(
        n4763) );
  AOI21_X1 U5310 ( .B1(n4764), .B2(keyinput_g92), .A(n4763), .ZN(n4783) );
  AOI22_X1 U5311 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_g42), .B1(
        D_REG_31__SCAN_IN), .B2(keyinput_g118), .ZN(n4765) );
  OAI221_X1 U5312 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_g42), .C1(
        D_REG_31__SCAN_IN), .C2(keyinput_g118), .A(n4765), .ZN(n4772) );
  AOI22_X1 U5313 ( .A1(IR_REG_30__SCAN_IN), .A2(keyinput_g85), .B1(
        D_REG_14__SCAN_IN), .B2(keyinput_g101), .ZN(n4766) );
  OAI221_X1 U5314 ( .B1(IR_REG_30__SCAN_IN), .B2(keyinput_g85), .C1(
        D_REG_14__SCAN_IN), .C2(keyinput_g101), .A(n4766), .ZN(n4771) );
  AOI22_X1 U5315 ( .A1(REG0_REG_3__SCAN_IN), .A2(keyinput_g122), .B1(
        IR_REG_31__SCAN_IN), .B2(keyinput_g86), .ZN(n4767) );
  OAI221_X1 U5316 ( .B1(REG0_REG_3__SCAN_IN), .B2(keyinput_g122), .C1(
        IR_REG_31__SCAN_IN), .C2(keyinput_g86), .A(n4767), .ZN(n4770) );
  AOI22_X1 U5317 ( .A1(REG0_REG_8__SCAN_IN), .A2(keyinput_g127), .B1(
        IR_REG_11__SCAN_IN), .B2(keyinput_g66), .ZN(n4768) );
  OAI221_X1 U5318 ( .B1(REG0_REG_8__SCAN_IN), .B2(keyinput_g127), .C1(
        IR_REG_11__SCAN_IN), .C2(keyinput_g66), .A(n4768), .ZN(n4769) );
  NOR4_X1 U5319 ( .A1(n4772), .A2(n4771), .A3(n4770), .A4(n4769), .ZN(n4782)
         );
  AOI22_X1 U5320 ( .A1(DATAI_6_), .A2(keyinput_g25), .B1(IR_REG_2__SCAN_IN), 
        .B2(keyinput_g57), .ZN(n4773) );
  OAI221_X1 U5321 ( .B1(DATAI_6_), .B2(keyinput_g25), .C1(IR_REG_2__SCAN_IN), 
        .C2(keyinput_g57), .A(n4773), .ZN(n4780) );
  AOI22_X1 U5322 ( .A1(DATAI_11_), .A2(keyinput_g20), .B1(D_REG_7__SCAN_IN), 
        .B2(keyinput_g94), .ZN(n4774) );
  OAI221_X1 U5323 ( .B1(DATAI_11_), .B2(keyinput_g20), .C1(D_REG_7__SCAN_IN), 
        .C2(keyinput_g94), .A(n4774), .ZN(n4779) );
  AOI22_X1 U5324 ( .A1(D_REG_4__SCAN_IN), .A2(keyinput_g91), .B1(
        D_REG_1__SCAN_IN), .B2(keyinput_g88), .ZN(n4775) );
  OAI221_X1 U5325 ( .B1(D_REG_4__SCAN_IN), .B2(keyinput_g91), .C1(
        D_REG_1__SCAN_IN), .C2(keyinput_g88), .A(n4775), .ZN(n4778) );
  AOI22_X1 U5326 ( .A1(REG3_REG_10__SCAN_IN), .A2(keyinput_g37), .B1(
        IR_REG_25__SCAN_IN), .B2(keyinput_g80), .ZN(n4776) );
  OAI221_X1 U5327 ( .B1(REG3_REG_10__SCAN_IN), .B2(keyinput_g37), .C1(
        IR_REG_25__SCAN_IN), .C2(keyinput_g80), .A(n4776), .ZN(n4777) );
  NOR4_X1 U5328 ( .A1(n4780), .A2(n4779), .A3(n4778), .A4(n4777), .ZN(n4781)
         );
  NAND4_X1 U5329 ( .A1(n4784), .A2(n4783), .A3(n4782), .A4(n4781), .ZN(n4898)
         );
  AOI22_X1 U5330 ( .A1(n5001), .A2(keyinput_g65), .B1(keyinput_g103), .B2(
        n4786), .ZN(n4785) );
  OAI221_X1 U5331 ( .B1(n5001), .B2(keyinput_g65), .C1(n4786), .C2(
        keyinput_g103), .A(n4785), .ZN(n4796) );
  INV_X1 U5332 ( .A(DATAI_4_), .ZN(n4789) );
  INV_X1 U5333 ( .A(DATAI_2_), .ZN(n4788) );
  AOI22_X1 U5334 ( .A1(n4789), .A2(keyinput_g27), .B1(n4788), .B2(keyinput_g29), .ZN(n4787) );
  OAI221_X1 U5335 ( .B1(n4789), .B2(keyinput_g27), .C1(n4788), .C2(
        keyinput_g29), .A(n4787), .ZN(n4795) );
  XOR2_X1 U5336 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_g41), .Z(n4792) );
  XNOR2_X1 U5337 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_g59), .ZN(n4791) );
  XNOR2_X1 U5338 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_g58), .ZN(n4790) );
  NAND3_X1 U5339 ( .A1(n4792), .A2(n4791), .A3(n4790), .ZN(n4794) );
  XNOR2_X1 U5340 ( .A(n5054), .B(keyinput_g116), .ZN(n4793) );
  NOR4_X1 U5341 ( .A1(n4796), .A2(n4795), .A3(n4794), .A4(n4793), .ZN(n4839)
         );
  XNOR2_X1 U5342 ( .A(n4797), .B(keyinput_g84), .ZN(n4803) );
  XNOR2_X1 U5343 ( .A(n4798), .B(keyinput_g62), .ZN(n4802) );
  XNOR2_X1 U5344 ( .A(n4799), .B(keyinput_g82), .ZN(n4801) );
  XNOR2_X1 U5345 ( .A(n4975), .B(keyinput_g49), .ZN(n4800) );
  NOR4_X1 U5346 ( .A1(n4803), .A2(n4802), .A3(n4801), .A4(n4800), .ZN(n4807)
         );
  XOR2_X1 U5347 ( .A(n5010), .B(keyinput_g125), .Z(n4806) );
  XNOR2_X1 U5348 ( .A(DATAI_3_), .B(keyinput_g28), .ZN(n4805) );
  XNOR2_X1 U5349 ( .A(IR_REG_17__SCAN_IN), .B(keyinput_g72), .ZN(n4804) );
  NAND4_X1 U5350 ( .A1(n4807), .A2(n4806), .A3(n4805), .A4(n4804), .ZN(n4810)
         );
  XNOR2_X1 U5351 ( .A(n4808), .B(keyinput_g99), .ZN(n4809) );
  NOR2_X1 U5352 ( .A1(n4810), .A2(n4809), .ZN(n4838) );
  AOI22_X1 U5353 ( .A1(n2487), .A2(keyinput_g77), .B1(keyinput_g112), .B2(
        n4812), .ZN(n4811) );
  OAI221_X1 U5354 ( .B1(n2487), .B2(keyinput_g77), .C1(n4812), .C2(
        keyinput_g112), .A(n4811), .ZN(n4823) );
  INV_X1 U5355 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4814) );
  AOI22_X1 U5356 ( .A1(n4815), .A2(keyinput_g98), .B1(keyinput_g34), .B2(n4814), .ZN(n4813) );
  OAI221_X1 U5357 ( .B1(n4815), .B2(keyinput_g98), .C1(n4814), .C2(
        keyinput_g34), .A(n4813), .ZN(n4822) );
  XNOR2_X1 U5358 ( .A(n5059), .B(keyinput_g102), .ZN(n4821) );
  XOR2_X1 U5359 ( .A(n4816), .B(keyinput_g19), .Z(n4819) );
  XNOR2_X1 U5360 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_g68), .ZN(n4818) );
  XNOR2_X1 U5361 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_g76), .ZN(n4817) );
  NAND3_X1 U5362 ( .A1(n4819), .A2(n4818), .A3(n4817), .ZN(n4820) );
  NOR4_X1 U5363 ( .A1(n4823), .A2(n4822), .A3(n4821), .A4(n4820), .ZN(n4837)
         );
  AOI22_X1 U5364 ( .A1(n5013), .A2(keyinput_g47), .B1(keyinput_g8), .B2(n4978), 
        .ZN(n4824) );
  OAI221_X1 U5365 ( .B1(n5013), .B2(keyinput_g47), .C1(n4978), .C2(keyinput_g8), .A(n4824), .ZN(n4835) );
  AOI22_X1 U5366 ( .A1(n4827), .A2(keyinput_g0), .B1(n4826), .B2(keyinput_g74), 
        .ZN(n4825) );
  OAI221_X1 U5367 ( .B1(n4827), .B2(keyinput_g0), .C1(n4826), .C2(keyinput_g74), .A(n4825), .ZN(n4834) );
  XOR2_X1 U5368 ( .A(n4828), .B(keyinput_g21), .Z(n4832) );
  XNOR2_X1 U5369 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_g60), .ZN(n4831) );
  XNOR2_X1 U5370 ( .A(DATAI_5_), .B(keyinput_g26), .ZN(n4830) );
  NAND4_X1 U5371 ( .A1(n4832), .A2(n4831), .A3(n4830), .A4(n4829), .ZN(n4833)
         );
  NOR3_X1 U5372 ( .A1(n4835), .A2(n4834), .A3(n4833), .ZN(n4836) );
  NAND4_X1 U5373 ( .A1(n4839), .A2(n4838), .A3(n4837), .A4(n4836), .ZN(n4897)
         );
  AOI22_X1 U5374 ( .A1(n4999), .A2(keyinput_g69), .B1(keyinput_g106), .B2(
        n4841), .ZN(n4840) );
  OAI221_X1 U5375 ( .B1(n4999), .B2(keyinput_g69), .C1(n4841), .C2(
        keyinput_g106), .A(n4840), .ZN(n4853) );
  INV_X1 U5376 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4844) );
  AOI22_X1 U5377 ( .A1(n4844), .A2(keyinput_g43), .B1(keyinput_g4), .B2(n4843), 
        .ZN(n4842) );
  OAI221_X1 U5378 ( .B1(n4844), .B2(keyinput_g43), .C1(n4843), .C2(keyinput_g4), .A(n4842), .ZN(n4852) );
  INV_X1 U5379 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4846) );
  AOI22_X1 U5380 ( .A1(n4847), .A2(keyinput_g97), .B1(keyinput_g40), .B2(n4846), .ZN(n4845) );
  OAI221_X1 U5381 ( .B1(n4847), .B2(keyinput_g97), .C1(n4846), .C2(
        keyinput_g40), .A(n4845), .ZN(n4851) );
  XOR2_X1 U5382 ( .A(n2790), .B(keyinput_g48), .Z(n4849) );
  XNOR2_X1 U5383 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_g50), .ZN(n4848) );
  NAND2_X1 U5384 ( .A1(n4849), .A2(n4848), .ZN(n4850) );
  NOR4_X1 U5385 ( .A1(n4853), .A2(n4852), .A3(n4851), .A4(n4850), .ZN(n4895)
         );
  AOI22_X1 U5386 ( .A1(n4856), .A2(keyinput_g119), .B1(n4855), .B2(
        keyinput_g117), .ZN(n4854) );
  OAI221_X1 U5387 ( .B1(n4856), .B2(keyinput_g119), .C1(n4855), .C2(
        keyinput_g117), .A(n4854), .ZN(n4864) );
  XOR2_X1 U5388 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_g63), .Z(n4863) );
  INV_X1 U5389 ( .A(IR_REG_16__SCAN_IN), .ZN(n4998) );
  XNOR2_X1 U5390 ( .A(keyinput_g71), .B(n4998), .ZN(n4862) );
  XNOR2_X1 U5391 ( .A(D_REG_0__SCAN_IN), .B(keyinput_g87), .ZN(n4860) );
  XNOR2_X1 U5392 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_g38), .ZN(n4859) );
  XNOR2_X1 U5393 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_g55), .ZN(n4858) );
  XNOR2_X1 U5394 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_g73), .ZN(n4857) );
  NAND4_X1 U5395 ( .A1(n4860), .A2(n4859), .A3(n4858), .A4(n4857), .ZN(n4861)
         );
  NOR4_X1 U5396 ( .A1(n4864), .A2(n4863), .A3(n4862), .A4(n4861), .ZN(n4894)
         );
  AOI22_X1 U5397 ( .A1(n4867), .A2(keyinput_g15), .B1(n4866), .B2(keyinput_g9), 
        .ZN(n4865) );
  OAI221_X1 U5398 ( .B1(n4867), .B2(keyinput_g15), .C1(n4866), .C2(keyinput_g9), .A(n4865), .ZN(n4877) );
  AOI22_X1 U5399 ( .A1(n5011), .A2(keyinput_g61), .B1(keyinput_g13), .B2(n4977), .ZN(n4868) );
  OAI221_X1 U5400 ( .B1(n5011), .B2(keyinput_g61), .C1(n4977), .C2(
        keyinput_g13), .A(n4868), .ZN(n4876) );
  AOI22_X1 U5401 ( .A1(n4871), .A2(keyinput_g108), .B1(keyinput_g51), .B2(
        n4870), .ZN(n4869) );
  OAI221_X1 U5402 ( .B1(n4871), .B2(keyinput_g108), .C1(n4870), .C2(
        keyinput_g51), .A(n4869), .ZN(n4875) );
  INV_X1 U5403 ( .A(DATAI_13_), .ZN(n4873) );
  AOI22_X1 U5404 ( .A1(n4873), .A2(keyinput_g18), .B1(n5038), .B2(keyinput_g95), .ZN(n4872) );
  OAI221_X1 U5405 ( .B1(n4873), .B2(keyinput_g18), .C1(n5038), .C2(
        keyinput_g95), .A(n4872), .ZN(n4874) );
  NOR4_X1 U5406 ( .A1(n4877), .A2(n4876), .A3(n4875), .A4(n4874), .ZN(n4893)
         );
  AOI22_X1 U5407 ( .A1(n4880), .A2(keyinput_g113), .B1(keyinput_g45), .B2(
        n4879), .ZN(n4878) );
  OAI221_X1 U5408 ( .B1(n4880), .B2(keyinput_g113), .C1(n4879), .C2(
        keyinput_g45), .A(n4878), .ZN(n4884) );
  XNOR2_X1 U5409 ( .A(n4881), .B(keyinput_g111), .ZN(n4883) );
  XOR2_X1 U5410 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_g64), .Z(n4882) );
  OR3_X1 U5411 ( .A1(n4884), .A2(n4883), .A3(n4882), .ZN(n4891) );
  INV_X1 U5412 ( .A(DATAI_29_), .ZN(n4887) );
  INV_X1 U5413 ( .A(DATAI_8_), .ZN(n4886) );
  AOI22_X1 U5414 ( .A1(n4887), .A2(keyinput_g2), .B1(keyinput_g23), .B2(n4886), 
        .ZN(n4885) );
  OAI221_X1 U5415 ( .B1(n4887), .B2(keyinput_g2), .C1(n4886), .C2(keyinput_g23), .A(n4885), .ZN(n4890) );
  AOI22_X1 U5416 ( .A1(n5061), .A2(keyinput_g121), .B1(n5069), .B2(
        keyinput_g39), .ZN(n4888) );
  OAI221_X1 U5417 ( .B1(n5061), .B2(keyinput_g121), .C1(n5069), .C2(
        keyinput_g39), .A(n4888), .ZN(n4889) );
  NOR3_X1 U5418 ( .A1(n4891), .A2(n4890), .A3(n4889), .ZN(n4892) );
  NAND4_X1 U5419 ( .A1(n4895), .A2(n4894), .A3(n4893), .A4(n4892), .ZN(n4896)
         );
  NOR4_X1 U5420 ( .A1(n4899), .A2(n4898), .A3(n4897), .A4(n4896), .ZN(n5096)
         );
  XOR2_X1 U5421 ( .A(keyinput_g115), .B(keyinput_f115), .Z(n5094) );
  XOR2_X1 U5422 ( .A(keyinput_f0), .B(DATAI_31_), .Z(n4906) );
  AOI22_X1 U5423 ( .A1(DATAI_25_), .A2(keyinput_f6), .B1(STATE_REG_SCAN_IN), 
        .B2(keyinput_f32), .ZN(n4900) );
  OAI221_X1 U5424 ( .B1(DATAI_25_), .B2(keyinput_f6), .C1(STATE_REG_SCAN_IN), 
        .C2(keyinput_f32), .A(n4900), .ZN(n4905) );
  AOI22_X1 U5425 ( .A1(DATAI_26_), .A2(keyinput_f5), .B1(DATAI_24_), .B2(
        keyinput_f7), .ZN(n4901) );
  OAI221_X1 U5426 ( .B1(DATAI_26_), .B2(keyinput_f5), .C1(DATAI_24_), .C2(
        keyinput_f7), .A(n4901), .ZN(n4904) );
  AOI22_X1 U5427 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput_f52), .B1(DATAI_19_), 
        .B2(keyinput_f12), .ZN(n4902) );
  OAI221_X1 U5428 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput_f52), .C1(DATAI_19_), .C2(keyinput_f12), .A(n4902), .ZN(n4903) );
  NOR4_X1 U5429 ( .A1(n4906), .A2(n4905), .A3(n4904), .A4(n4903), .ZN(n4934)
         );
  AOI22_X1 U5430 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput_f34), .B1(
        REG3_REG_28__SCAN_IN), .B2(keyinput_f40), .ZN(n4907) );
  OAI221_X1 U5431 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput_f34), .C1(
        REG3_REG_28__SCAN_IN), .C2(keyinput_f40), .A(n4907), .ZN(n4914) );
  AOI22_X1 U5432 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(REG3_REG_20__SCAN_IN), 
        .B2(keyinput_f53), .ZN(n4908) );
  OAI221_X1 U5433 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(REG3_REG_20__SCAN_IN), .C2(keyinput_f53), .A(n4908), .ZN(n4913) );
  AOI22_X1 U5434 ( .A1(DATAI_22_), .A2(keyinput_f9), .B1(DATAI_27_), .B2(
        keyinput_f4), .ZN(n4909) );
  OAI221_X1 U5435 ( .B1(DATAI_22_), .B2(keyinput_f9), .C1(DATAI_27_), .C2(
        keyinput_f4), .A(n4909), .ZN(n4912) );
  AOI22_X1 U5436 ( .A1(DATAI_20_), .A2(keyinput_f11), .B1(DATAI_21_), .B2(
        keyinput_f10), .ZN(n4910) );
  OAI221_X1 U5437 ( .B1(DATAI_20_), .B2(keyinput_f11), .C1(DATAI_21_), .C2(
        keyinput_f10), .A(n4910), .ZN(n4911) );
  NOR4_X1 U5438 ( .A1(n4914), .A2(n4913), .A3(n4912), .A4(n4911), .ZN(n4933)
         );
  AOI22_X1 U5439 ( .A1(DATAI_17_), .A2(keyinput_f14), .B1(REG3_REG_7__SCAN_IN), 
        .B2(keyinput_f33), .ZN(n4915) );
  OAI221_X1 U5440 ( .B1(DATAI_17_), .B2(keyinput_f14), .C1(REG3_REG_7__SCAN_IN), .C2(keyinput_f33), .A(n4915), .ZN(n4922) );
  AOI22_X1 U5441 ( .A1(REG3_REG_14__SCAN_IN), .A2(keyinput_f35), .B1(
        D_REG_31__SCAN_IN), .B2(keyinput_f118), .ZN(n4916) );
  OAI221_X1 U5442 ( .B1(REG3_REG_14__SCAN_IN), .B2(keyinput_f35), .C1(
        D_REG_31__SCAN_IN), .C2(keyinput_f118), .A(n4916), .ZN(n4921) );
  AOI22_X1 U5443 ( .A1(D_REG_14__SCAN_IN), .A2(keyinput_f101), .B1(
        D_REG_27__SCAN_IN), .B2(keyinput_f114), .ZN(n4917) );
  OAI221_X1 U5444 ( .B1(D_REG_14__SCAN_IN), .B2(keyinput_f101), .C1(
        D_REG_27__SCAN_IN), .C2(keyinput_f114), .A(n4917), .ZN(n4920) );
  AOI22_X1 U5445 ( .A1(D_REG_2__SCAN_IN), .A2(keyinput_f89), .B1(
        D_REG_13__SCAN_IN), .B2(keyinput_f100), .ZN(n4918) );
  OAI221_X1 U5446 ( .B1(D_REG_2__SCAN_IN), .B2(keyinput_f89), .C1(
        D_REG_13__SCAN_IN), .C2(keyinput_f100), .A(n4918), .ZN(n4919) );
  NOR4_X1 U5447 ( .A1(n4922), .A2(n4921), .A3(n4920), .A4(n4919), .ZN(n4932)
         );
  AOI22_X1 U5448 ( .A1(REG0_REG_3__SCAN_IN), .A2(keyinput_f122), .B1(DATAI_7_), 
        .B2(keyinput_f24), .ZN(n4923) );
  OAI221_X1 U5449 ( .B1(REG0_REG_3__SCAN_IN), .B2(keyinput_f122), .C1(DATAI_7_), .C2(keyinput_f24), .A(n4923), .ZN(n4930) );
  AOI22_X1 U5450 ( .A1(REG0_REG_4__SCAN_IN), .A2(keyinput_f123), .B1(
        REG0_REG_5__SCAN_IN), .B2(keyinput_f124), .ZN(n4924) );
  OAI221_X1 U5451 ( .B1(REG0_REG_4__SCAN_IN), .B2(keyinput_f123), .C1(
        REG0_REG_5__SCAN_IN), .C2(keyinput_f124), .A(n4924), .ZN(n4929) );
  AOI22_X1 U5452 ( .A1(REG0_REG_7__SCAN_IN), .A2(keyinput_f126), .B1(
        REG0_REG_8__SCAN_IN), .B2(keyinput_f127), .ZN(n4925) );
  OAI221_X1 U5453 ( .B1(REG0_REG_7__SCAN_IN), .B2(keyinput_f126), .C1(
        REG0_REG_8__SCAN_IN), .C2(keyinput_f127), .A(n4925), .ZN(n4928) );
  AOI22_X1 U5454 ( .A1(DATAI_12_), .A2(keyinput_f19), .B1(IR_REG_28__SCAN_IN), 
        .B2(keyinput_f83), .ZN(n4926) );
  OAI221_X1 U5455 ( .B1(DATAI_12_), .B2(keyinput_f19), .C1(IR_REG_28__SCAN_IN), 
        .C2(keyinput_f83), .A(n4926), .ZN(n4927) );
  NOR4_X1 U5456 ( .A1(n4930), .A2(n4929), .A3(n4928), .A4(n4927), .ZN(n4931)
         );
  NAND4_X1 U5457 ( .A1(n4934), .A2(n4933), .A3(n4932), .A4(n4931), .ZN(n5090)
         );
  AOI22_X1 U5458 ( .A1(IR_REG_11__SCAN_IN), .A2(keyinput_f66), .B1(
        IR_REG_13__SCAN_IN), .B2(keyinput_f68), .ZN(n4935) );
  OAI221_X1 U5459 ( .B1(IR_REG_11__SCAN_IN), .B2(keyinput_f66), .C1(
        IR_REG_13__SCAN_IN), .C2(keyinput_f68), .A(n4935), .ZN(n4942) );
  AOI22_X1 U5460 ( .A1(DATAI_5_), .A2(keyinput_f26), .B1(DATAI_10_), .B2(
        keyinput_f21), .ZN(n4936) );
  OAI221_X1 U5461 ( .B1(DATAI_5_), .B2(keyinput_f26), .C1(DATAI_10_), .C2(
        keyinput_f21), .A(n4936), .ZN(n4941) );
  AOI22_X1 U5462 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput_f50), .B1(
        IR_REG_3__SCAN_IN), .B2(keyinput_f58), .ZN(n4937) );
  OAI221_X1 U5463 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput_f50), .C1(
        IR_REG_3__SCAN_IN), .C2(keyinput_f58), .A(n4937), .ZN(n4940) );
  AOI22_X1 U5464 ( .A1(REG0_REG_0__SCAN_IN), .A2(keyinput_f119), .B1(
        IR_REG_2__SCAN_IN), .B2(keyinput_f57), .ZN(n4938) );
  OAI221_X1 U5465 ( .B1(REG0_REG_0__SCAN_IN), .B2(keyinput_f119), .C1(
        IR_REG_2__SCAN_IN), .C2(keyinput_f57), .A(n4938), .ZN(n4939) );
  NOR4_X1 U5466 ( .A1(n4942), .A2(n4941), .A3(n4940), .A4(n4939), .ZN(n4970)
         );
  AOI22_X1 U5467 ( .A1(DATAI_8_), .A2(keyinput_f23), .B1(IR_REG_8__SCAN_IN), 
        .B2(keyinput_f63), .ZN(n4943) );
  OAI221_X1 U5468 ( .B1(DATAI_8_), .B2(keyinput_f23), .C1(IR_REG_8__SCAN_IN), 
        .C2(keyinput_f63), .A(n4943), .ZN(n4950) );
  AOI22_X1 U5469 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput_f51), .B1(
        IR_REG_9__SCAN_IN), .B2(keyinput_f64), .ZN(n4944) );
  OAI221_X1 U5470 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput_f51), .C1(
        IR_REG_9__SCAN_IN), .C2(keyinput_f64), .A(n4944), .ZN(n4949) );
  AOI22_X1 U5471 ( .A1(D_REG_19__SCAN_IN), .A2(keyinput_f106), .B1(
        IR_REG_20__SCAN_IN), .B2(keyinput_f75), .ZN(n4945) );
  OAI221_X1 U5472 ( .B1(D_REG_19__SCAN_IN), .B2(keyinput_f106), .C1(
        IR_REG_20__SCAN_IN), .C2(keyinput_f75), .A(n4945), .ZN(n4948) );
  AOI22_X1 U5473 ( .A1(D_REG_12__SCAN_IN), .A2(keyinput_f99), .B1(
        D_REG_25__SCAN_IN), .B2(keyinput_f112), .ZN(n4946) );
  OAI221_X1 U5474 ( .B1(D_REG_12__SCAN_IN), .B2(keyinput_f99), .C1(
        D_REG_25__SCAN_IN), .C2(keyinput_f112), .A(n4946), .ZN(n4947) );
  NOR4_X1 U5475 ( .A1(n4950), .A2(n4949), .A3(n4948), .A4(n4947), .ZN(n4969)
         );
  AOI22_X1 U5476 ( .A1(D_REG_10__SCAN_IN), .A2(keyinput_f97), .B1(
        D_REG_5__SCAN_IN), .B2(keyinput_f92), .ZN(n4951) );
  OAI221_X1 U5477 ( .B1(D_REG_10__SCAN_IN), .B2(keyinput_f97), .C1(
        D_REG_5__SCAN_IN), .C2(keyinput_f92), .A(n4951), .ZN(n4958) );
  AOI22_X1 U5478 ( .A1(D_REG_16__SCAN_IN), .A2(keyinput_f103), .B1(
        D_REG_11__SCAN_IN), .B2(keyinput_f98), .ZN(n4952) );
  OAI221_X1 U5479 ( .B1(D_REG_16__SCAN_IN), .B2(keyinput_f103), .C1(
        D_REG_11__SCAN_IN), .C2(keyinput_f98), .A(n4952), .ZN(n4957) );
  AOI22_X1 U5480 ( .A1(D_REG_21__SCAN_IN), .A2(keyinput_f108), .B1(
        D_REG_30__SCAN_IN), .B2(keyinput_f117), .ZN(n4953) );
  OAI221_X1 U5481 ( .B1(D_REG_21__SCAN_IN), .B2(keyinput_f108), .C1(
        D_REG_30__SCAN_IN), .C2(keyinput_f117), .A(n4953), .ZN(n4956) );
  AOI22_X1 U5482 ( .A1(D_REG_26__SCAN_IN), .A2(keyinput_f113), .B1(
        D_REG_24__SCAN_IN), .B2(keyinput_f111), .ZN(n4954) );
  OAI221_X1 U5483 ( .B1(D_REG_26__SCAN_IN), .B2(keyinput_f113), .C1(
        D_REG_24__SCAN_IN), .C2(keyinput_f111), .A(n4954), .ZN(n4955) );
  NOR4_X1 U5484 ( .A1(n4958), .A2(n4957), .A3(n4956), .A4(n4955), .ZN(n4968)
         );
  AOI22_X1 U5485 ( .A1(REG3_REG_17__SCAN_IN), .A2(keyinput_f48), .B1(
        REG3_REG_25__SCAN_IN), .B2(keyinput_f45), .ZN(n4959) );
  OAI221_X1 U5486 ( .B1(REG3_REG_17__SCAN_IN), .B2(keyinput_f48), .C1(
        REG3_REG_25__SCAN_IN), .C2(keyinput_f45), .A(n4959), .ZN(n4966) );
  AOI22_X1 U5487 ( .A1(REG3_REG_8__SCAN_IN), .A2(keyinput_f41), .B1(
        REG3_REG_12__SCAN_IN), .B2(keyinput_f44), .ZN(n4960) );
  OAI221_X1 U5488 ( .B1(REG3_REG_8__SCAN_IN), .B2(keyinput_f41), .C1(
        REG3_REG_12__SCAN_IN), .C2(keyinput_f44), .A(n4960), .ZN(n4965) );
  AOI22_X1 U5489 ( .A1(DATAI_16_), .A2(keyinput_f15), .B1(IR_REG_26__SCAN_IN), 
        .B2(keyinput_f81), .ZN(n4961) );
  OAI221_X1 U5490 ( .B1(DATAI_16_), .B2(keyinput_f15), .C1(IR_REG_26__SCAN_IN), 
        .C2(keyinput_f81), .A(n4961), .ZN(n4964) );
  AOI22_X1 U5491 ( .A1(DATAI_13_), .A2(keyinput_f18), .B1(DATAI_29_), .B2(
        keyinput_f2), .ZN(n4962) );
  OAI221_X1 U5492 ( .B1(DATAI_13_), .B2(keyinput_f18), .C1(DATAI_29_), .C2(
        keyinput_f2), .A(n4962), .ZN(n4963) );
  NOR4_X1 U5493 ( .A1(n4966), .A2(n4965), .A3(n4964), .A4(n4963), .ZN(n4967)
         );
  NAND4_X1 U5494 ( .A1(n4970), .A2(n4969), .A3(n4968), .A4(n4967), .ZN(n5089)
         );
  AOI22_X1 U5495 ( .A1(REG3_REG_21__SCAN_IN), .A2(keyinput_f43), .B1(
        IR_REG_25__SCAN_IN), .B2(keyinput_f80), .ZN(n4971) );
  OAI221_X1 U5496 ( .B1(REG3_REG_21__SCAN_IN), .B2(keyinput_f43), .C1(
        IR_REG_25__SCAN_IN), .C2(keyinput_f80), .A(n4971), .ZN(n4982) );
  AOI22_X1 U5497 ( .A1(DATAI_4_), .A2(keyinput_f27), .B1(IR_REG_23__SCAN_IN), 
        .B2(keyinput_f78), .ZN(n4972) );
  OAI221_X1 U5498 ( .B1(DATAI_4_), .B2(keyinput_f27), .C1(IR_REG_23__SCAN_IN), 
        .C2(keyinput_f78), .A(n4972), .ZN(n4981) );
  AOI22_X1 U5499 ( .A1(n4975), .A2(keyinput_f49), .B1(keyinput_f3), .B2(n4974), 
        .ZN(n4973) );
  OAI221_X1 U5500 ( .B1(n4975), .B2(keyinput_f49), .C1(n4974), .C2(keyinput_f3), .A(n4973), .ZN(n4980) );
  AOI22_X1 U5501 ( .A1(n4978), .A2(keyinput_f8), .B1(keyinput_f13), .B2(n4977), 
        .ZN(n4976) );
  OAI221_X1 U5502 ( .B1(n4978), .B2(keyinput_f8), .C1(n4977), .C2(keyinput_f13), .A(n4976), .ZN(n4979) );
  NOR4_X1 U5503 ( .A1(n4982), .A2(n4981), .A3(n4980), .A4(n4979), .ZN(n5025)
         );
  XOR2_X1 U5504 ( .A(n3247), .B(keyinput_f42), .Z(n4987) );
  XOR2_X1 U5505 ( .A(n4983), .B(keyinput_f16), .Z(n4986) );
  XNOR2_X1 U5506 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_f86), .ZN(n4985) );
  XNOR2_X1 U5507 ( .A(IR_REG_30__SCAN_IN), .B(keyinput_f85), .ZN(n4984) );
  NAND4_X1 U5508 ( .A1(n4987), .A2(n4986), .A3(n4985), .A4(n4984), .ZN(n4993)
         );
  XNOR2_X1 U5509 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput_f54), .ZN(n4991) );
  XNOR2_X1 U5510 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_f38), .ZN(n4990) );
  XNOR2_X1 U5511 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_f82), .ZN(n4989) );
  XNOR2_X1 U5512 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_f55), .ZN(n4988) );
  NAND4_X1 U5513 ( .A1(n4991), .A2(n4990), .A3(n4989), .A4(n4988), .ZN(n4992)
         );
  NOR2_X1 U5514 ( .A1(n4993), .A2(n4992), .ZN(n5024) );
  AOI22_X1 U5515 ( .A1(n4996), .A2(keyinput_f70), .B1(keyinput_f17), .B2(n4995), .ZN(n4994) );
  OAI221_X1 U5516 ( .B1(n4996), .B2(keyinput_f70), .C1(n4995), .C2(
        keyinput_f17), .A(n4994), .ZN(n5008) );
  AOI22_X1 U5517 ( .A1(n4999), .A2(keyinput_f69), .B1(n4998), .B2(keyinput_f71), .ZN(n4997) );
  OAI221_X1 U5518 ( .B1(n4999), .B2(keyinput_f69), .C1(n4998), .C2(
        keyinput_f71), .A(n4997), .ZN(n5007) );
  INV_X1 U5519 ( .A(IR_REG_12__SCAN_IN), .ZN(n5002) );
  AOI22_X1 U5520 ( .A1(n5002), .A2(keyinput_f67), .B1(keyinput_f65), .B2(n5001), .ZN(n5000) );
  OAI221_X1 U5521 ( .B1(n5002), .B2(keyinput_f67), .C1(n5001), .C2(
        keyinput_f65), .A(n5000), .ZN(n5006) );
  XNOR2_X1 U5522 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_f73), .ZN(n5004) );
  XNOR2_X1 U5523 ( .A(IR_REG_17__SCAN_IN), .B(keyinput_f72), .ZN(n5003) );
  NAND2_X1 U5524 ( .A1(n5004), .A2(n5003), .ZN(n5005) );
  NOR4_X1 U5525 ( .A1(n5008), .A2(n5007), .A3(n5006), .A4(n5005), .ZN(n5023)
         );
  AOI22_X1 U5526 ( .A1(n5011), .A2(keyinput_f61), .B1(keyinput_f125), .B2(
        n5010), .ZN(n5009) );
  OAI221_X1 U5527 ( .B1(n5011), .B2(keyinput_f61), .C1(n5010), .C2(
        keyinput_f125), .A(n5009), .ZN(n5021) );
  INV_X1 U5528 ( .A(DATAI_6_), .ZN(n5012) );
  XNOR2_X1 U5529 ( .A(keyinput_f25), .B(n5012), .ZN(n5020) );
  XNOR2_X1 U5530 ( .A(keyinput_f47), .B(n5013), .ZN(n5019) );
  XNOR2_X1 U5531 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_f60), .ZN(n5017) );
  XNOR2_X1 U5532 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_f62), .ZN(n5016) );
  XNOR2_X1 U5533 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_f59), .ZN(n5015) );
  XNOR2_X1 U5534 ( .A(DATAI_0_), .B(keyinput_f31), .ZN(n5014) );
  NAND4_X1 U5535 ( .A1(n5017), .A2(n5016), .A3(n5015), .A4(n5014), .ZN(n5018)
         );
  NOR4_X1 U5536 ( .A1(n5021), .A2(n5020), .A3(n5019), .A4(n5018), .ZN(n5022)
         );
  NAND4_X1 U5537 ( .A1(n5025), .A2(n5024), .A3(n5023), .A4(n5022), .ZN(n5088)
         );
  XOR2_X1 U5538 ( .A(n5026), .B(keyinput_f120), .Z(n5030) );
  XNOR2_X1 U5539 ( .A(keyinput_f29), .B(DATAI_2_), .ZN(n5029) );
  XNOR2_X1 U5540 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_f76), .ZN(n5028) );
  XNOR2_X1 U5541 ( .A(IR_REG_19__SCAN_IN), .B(keyinput_f74), .ZN(n5027) );
  NAND4_X1 U5542 ( .A1(n5030), .A2(n5029), .A3(n5028), .A4(n5027), .ZN(n5036)
         );
  XNOR2_X1 U5543 ( .A(DATAI_1_), .B(keyinput_f30), .ZN(n5033) );
  XNOR2_X1 U5544 ( .A(DATAI_3_), .B(keyinput_f28), .ZN(n5032) );
  XNOR2_X1 U5545 ( .A(DATAI_11_), .B(keyinput_f20), .ZN(n5031) );
  NAND4_X1 U5546 ( .A1(n5034), .A2(n5033), .A3(n5032), .A4(n5031), .ZN(n5035)
         );
  NOR2_X1 U5547 ( .A1(n5036), .A2(n5035), .ZN(n5086) );
  AOI22_X1 U5548 ( .A1(n2487), .A2(keyinput_f77), .B1(keyinput_f95), .B2(n5038), .ZN(n5037) );
  OAI221_X1 U5549 ( .B1(n2487), .B2(keyinput_f77), .C1(n5038), .C2(
        keyinput_f95), .A(n5037), .ZN(n5051) );
  AOI22_X1 U5550 ( .A1(n5041), .A2(keyinput_f96), .B1(keyinput_f105), .B2(
        n5040), .ZN(n5039) );
  OAI221_X1 U5551 ( .B1(n5041), .B2(keyinput_f96), .C1(n5040), .C2(
        keyinput_f105), .A(n5039), .ZN(n5050) );
  AOI22_X1 U5552 ( .A1(n5044), .A2(keyinput_f104), .B1(keyinput_f109), .B2(
        n5043), .ZN(n5042) );
  OAI221_X1 U5553 ( .B1(n5044), .B2(keyinput_f104), .C1(n5043), .C2(
        keyinput_f109), .A(n5042), .ZN(n5049) );
  AOI22_X1 U5554 ( .A1(n5047), .A2(keyinput_f107), .B1(keyinput_f110), .B2(
        n5046), .ZN(n5045) );
  OAI221_X1 U5555 ( .B1(n5047), .B2(keyinput_f107), .C1(n5046), .C2(
        keyinput_f110), .A(n5045), .ZN(n5048) );
  NOR4_X1 U5556 ( .A1(n5051), .A2(n5050), .A3(n5049), .A4(n5048), .ZN(n5085)
         );
  AOI22_X1 U5557 ( .A1(n5054), .A2(keyinput_f116), .B1(keyinput_f93), .B2(
        n5053), .ZN(n5052) );
  OAI221_X1 U5558 ( .B1(n5054), .B2(keyinput_f116), .C1(n5053), .C2(
        keyinput_f93), .A(n5052), .ZN(n5067) );
  AOI22_X1 U5559 ( .A1(n5057), .A2(keyinput_f90), .B1(keyinput_f94), .B2(n5056), .ZN(n5055) );
  OAI221_X1 U5560 ( .B1(n5057), .B2(keyinput_f90), .C1(n5056), .C2(
        keyinput_f94), .A(n5055), .ZN(n5066) );
  AOI22_X1 U5561 ( .A1(n5060), .A2(keyinput_f91), .B1(n5059), .B2(
        keyinput_f102), .ZN(n5058) );
  OAI221_X1 U5562 ( .B1(n5060), .B2(keyinput_f91), .C1(n5059), .C2(
        keyinput_f102), .A(n5058), .ZN(n5065) );
  XOR2_X1 U5563 ( .A(n5061), .B(keyinput_f121), .Z(n5063) );
  XNOR2_X1 U5564 ( .A(IR_REG_29__SCAN_IN), .B(keyinput_f84), .ZN(n5062) );
  NAND2_X1 U5565 ( .A1(n5063), .A2(n5062), .ZN(n5064) );
  NOR4_X1 U5566 ( .A1(n5067), .A2(n5066), .A3(n5065), .A4(n5064), .ZN(n5084)
         );
  AOI22_X1 U5567 ( .A1(n5070), .A2(keyinput_f88), .B1(keyinput_f39), .B2(n5069), .ZN(n5068) );
  OAI221_X1 U5568 ( .B1(n5070), .B2(keyinput_f88), .C1(n5069), .C2(
        keyinput_f39), .A(n5068), .ZN(n5082) );
  AOI22_X1 U5569 ( .A1(n5073), .A2(keyinput_f46), .B1(n5072), .B2(keyinput_f36), .ZN(n5071) );
  OAI221_X1 U5570 ( .B1(n5073), .B2(keyinput_f46), .C1(n5072), .C2(
        keyinput_f36), .A(n5071), .ZN(n5081) );
  AOI22_X1 U5571 ( .A1(n2394), .A2(keyinput_f79), .B1(keyinput_f87), .B2(n5075), .ZN(n5074) );
  OAI221_X1 U5572 ( .B1(n2394), .B2(keyinput_f79), .C1(n5075), .C2(
        keyinput_f87), .A(n5074), .ZN(n5080) );
  INV_X1 U5573 ( .A(DATAI_9_), .ZN(n5078) );
  INV_X1 U5574 ( .A(REG3_REG_10__SCAN_IN), .ZN(n5077) );
  AOI22_X1 U5575 ( .A1(n5078), .A2(keyinput_f22), .B1(n5077), .B2(keyinput_f37), .ZN(n5076) );
  OAI221_X1 U5576 ( .B1(n5078), .B2(keyinput_f22), .C1(n5077), .C2(
        keyinput_f37), .A(n5076), .ZN(n5079) );
  NOR4_X1 U5577 ( .A1(n5082), .A2(n5081), .A3(n5080), .A4(n5079), .ZN(n5083)
         );
  NAND4_X1 U5578 ( .A1(n5086), .A2(n5085), .A3(n5084), .A4(n5083), .ZN(n5087)
         );
  NOR4_X1 U5579 ( .A1(n5090), .A2(n5089), .A3(n5088), .A4(n5087), .ZN(n5093)
         );
  NAND2_X1 U5580 ( .A1(keyinput_g115), .A2(n5092), .ZN(n5091) );
  OAI221_X1 U5581 ( .B1(n5094), .B2(n5093), .C1(keyinput_g115), .C2(n5092), 
        .A(n5091), .ZN(n5095) );
  AOI21_X1 U5582 ( .B1(n5097), .B2(n5096), .A(n5095), .ZN(n5099) );
  AOI22_X1 U5583 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n5098) );
  XNOR2_X1 U5584 ( .A(n5099), .B(n5098), .ZN(U3352) );
  CLKBUF_X1 U2481 ( .A(n2948), .Z(n2233) );
  CLKBUF_X1 U2482 ( .A(n2546), .Z(n3895) );
  CLKBUF_X1 U4847 ( .A(n4193), .Z(n4194) );
endmodule

